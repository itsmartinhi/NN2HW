library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
    port (
        in_rom_input_index:     in std_logic_vector(7 downto 0); -- the given rom input index
        in_rom_neuron_index:    in std_logic_vector(3 downto 0); -- the given neuron index
        out_data_rom:           out std_logic_vector(31 downto 0) -- the output datastream
    );
end ROM;

architecture RTL of ROM is 
    type t_rom_arr is array (0 to 2500) of std_logic_vector (31 downto 0);
    constant rom_arr: t_rom_arr := (
        -- here follows the generated array allocation
		"01010000000000000000000000000000",
		"01110110011101000111001001111000",
		"01111000011101010111011001110001",
		"01110100011110000111001101110010",
		"01110101011100110111011001110101",
		"01110001011110010111100001110110",
		"01111001011100010111010101110111",
		"01110101011101100111100101110010",
		"01111000011101110111010101110110",
		"01110110011101100111001101110010",
		"01110101011100010111011101111001",
		"01110100011100000111100001111001",
		"01111000011110010111101001111100",
		"01110001011100010111011101110111",
		"01110010011110010111010001110101",
		"01111001011101010111100001110010",
		"01110101011100010111100001111000",
		"01110011011100100111010101110101",
		"01100111011010110110111001110110",
		"01110001011100000110110101101100",
		"01110011011100100111000101101110",
		"01110001011101010111010101111001",
		"01111000011100100111011101110010",
		"01100111011011010110111001111001",
		"01111100011110110111010001110101",
		"10000011100100011000111101111010",
		"01110010011101101000101010001111",
		"01110011011011010110100101110010",
		"01110001011101000111011101110100",
		"01110111011100010111100001110001",
		"01110110011001110110101001110010",
		"10100000011111111000011001111000",
		"10011000100001011001011010001001",
		"10000001100010111001011110000111",
		"01110101011110100111010001111001",
		"01111001011101000111000101101100",
		"01110101011101100111011101110111",
		"01111011011101010110010101110101",
		"10010011100110011000010010000001",
		"10000001100100001001000101110100",
		"10001001100101011001001110000101",
		"01101100011110101000000001110010",
		"01110010011100000110011101100110",
		"01111000011101110111001101110110",
		"01111110100000010111000001101111",
		"01110111011111000110100001111111",
		"01110010100011111001000001101111",
		"01111101100011101000000010001101",
		"01110011100111111001100110001000",
		"01110110011011000101110001011110",
		"01110100011110000111001001110011",
		"10000111100000110111011101110001",
		"10001000100000101000100001110000",
		"01110011011111001000011001110100",
		"10001000100100101001010101110000",
		"10010001011100110111110001111000",
		"01110001011001000101110101110001",
		"01110111011100010111010101111001",
		"01111010011110100111010101101100",
		"01110100011110101000111110000001",
		"10001101100011100110111010001100",
		"01110111100001111000111110101100",
		"10101000100011001001000010010000",
		"01110111011001100101011010001111",
		"01111110011100100111100101110011",
		"01110101011100010111011101110001",
		"01110010100100100111110101110000",
		"01100010011101011001111101110010",
		"10011001100100111001000010001000",
		"10011011011100110111011110001110",
		"01110010011001110101111110100011",
		"01111001011101110111000101110010",
		"01111100011110011000011101110011",
		"10001101011100111001001001111001",
		"01101110100011111000110101111001",
		"01110011100101101011011001111111",
		"10011000100101001000100110001110",
		"01110110011001010110000110100000",
		"01110101011101100111001101111000",
		"10010000100001110110111001101101",
		"10001000011111110111001010001111",
		"01011011011011001000001001101000",
		"10000010011010010111001101011100",
		"10001101100101001010000110001111",
		"01110100011001110110011110010010",
		"01110100011101000111010001111001",
		"10001110101000010111011101110000",
		"10000100100000110111111001111111",
		"01011001011000011000011010101000",
		"10001101011101000111001101011110",
		"10010011100101001001000110010000",
		"01111000011011100111000110101110",
		"01110101011100110111101001110001",
		"10010110100111010111100110000100",
		"01111010100111010111111110001001",
		"01010011010110010110011010000010",
		"01111001011110010110111001011011",
		"10010111100011010111110101101001",
		"01110110011100011000000110011011",
		"01101010011100100111011101110110",
		"10100001100010001001001001110000",
		"10011110011011101000111010000110",
		"01011001010110000110110110101111",
		"01110100011110000111000101011001",
		"10011000100000111000111010000111",
		"01111001011101111000010010100000",
		"01100111011100000111100101110110",
		"10011101011101001001100110001010",
		"01101100100111111001000010010010",
		"01011010010011100110010001110011",
		"01110011011111100111000001100010",
		"10010010100010001000001110010001",
		"01110110011100000111110010011001",
		"01110010011100110111100001110100",
		"10001111100100001001010010001000",
		"10010111100011001001000110011001",
		"01101010010111000101100001101011",
		"10000000100000101000001001101011",
		"10001000100011001000100110010001",
		"01110010011101000110101110000010",
		"01110101011101000111100101110010",
		"10001111100110011001000110000101",
		"10000010101100001001011101111001",
		"01101000011000100101111001110100",
		"10000000011101001001110101110010",
		"10000011100010110111100110001101",
		"01110101011100010110111101111101",
		"01110000011101010111100101111000",
		"10000101100011000111111110000001",
		"01111010101001111001011110011001",
		"01110000011010000110000001101110",
		"01110001011101010111101001110101",
		"10000011100100100111010101101111",
		"01110011011110000111000001111011",
		"01101101011100010111011001110010",
		"10010010100100111000001101111110",
		"10011100100011010111101110010010",
		"01101101011011000110100010011010",
		"01101110100000110111111101101001",
		"01111110100110011000110110000001",
		"01111001011100110111000101110111",
		"01101111011110010111010101110110",
		"10001010100100001001010010000011",
		"10010011100101111001001110010100",
		"10000000011100101000100010100111",
		"10000000011111101000000101101101",
		"01101101100101011000100001111111",
		"01110101011101000111001001101110",
		"01110110011100010111011001110110",
		"10010011100011001000011001110101",
		"10001101100010100111110101111000",
		"01111011011100000111010010010011",
		"01110010011100110110111001111100",
		"01101110011111110111101101111001",
		"01110100011111010111001001101000",
		"01110110011101010111011101110111",
		"01111111100011001000000001011110",
		"01110111100010101000100110001100",
		"10000001011110011010100110000010",
		"10000101011100111000101101111110",
		"01110111100001000111011001111001",
		"01110100011100010110111101101000",
		"01110011011110010111011001110011",
		"10001101011110000110100001100000",
		"10011001100110011000111110000101",
		"01111110100010011000011110000101",
		"01101110011100001000111001110010",
		"01101110011101000110100101100110",
		"01110001011100100111010001101101",
		"01110101011101000111100001110101",
		"01101100011011100111001001110010",
		"01110101100011001000011101111011",
		"10001101100110001001101110011110",
		"01100000011101001000001110000011",
		"01110100011010000110010101011011",
		"01110101011101100111001101110001",
		"01110111011101000111011101111001",
		"01101010011011000110111101110000",
		"01100010010111010110011101100110",
		"01011011010110110110000101011110",
		"01100101010110110101101101100100",
		"01110111011011010110011001100110",
		"01110001011110000111100001111000",
		"01110110011100010111011101110100",
		"01110101011101100111011001110001",
		"01110100011011100111000001101111",
		"01101110011011100110101101110110",
		"01110000011100010110110001101110",
		"01110111011100010110110001101110",
		"01110111011101000111100101111001",
		"01110111011101010111100101110001",
		"01110100011110010111010001111001",
		"01110100011100100111011101110011",
		"01110011011100010111100101110001",
		"01111001011110000111011001110101",
		"01110101011011010111011001110101",
		"01110001011101010111100001111010",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"10111001000000000000000000000000",
		"01111000011101000111010001110111",
		"01110010011110010111001001110011",
		"01110110011100010111000101110100",
		"01111000011101110111000101110001",
		"01111000011101110111000101110111",
		"01110100011100010111011101110111",
		"01110110011110010111010001110111",
		"01110111011101000111100001110011",
		"01110010011101110111010101111000",
		"01111010011110000111011001110100",
		"01111010011110100111011101110001",
		"01111010011101010111001101110100",
		"01110101011101000111000101111001",
		"01111001011100100111001101110001",
		"01110110011101100111100101111000",
		"01110100011100100111100001110100",
		"01110000011011010110111101110101",
		"10010010011111111000001101110001",
		"01110100011110000111011010001000",
		"01111001011100110111000101111000",
		"01111001011110000111100101110101",
		"01110111011100000111011001110011",
		"01110100011101000111100001110100",
		"01100010011001100110111001110000",
		"10000100011101000111110001110101",
		"01110100011001110111011010001101",
		"01101111011011010110101001110010",
		"01110011011101010111011101110000",
		"01110010011101110111100001110100",
		"01110010011111100111101001110001",
		"01110110011110010111001101111100",
		"10000111100010101001000110000011",
		"10000011011111001000001110001010",
		"01101010011011010111100101111110",
		"01110110011100110110100101010101",
		"01111010011110000111001001110111",
		"01111001100001001000000001111010",
		"01101010011100010110100001100111",
		"10000101011101010111101001101101",
		"01111101011111010110101001111100",
		"01111111100010101000100001111111",
		"01110111011011110110001101101110",
		"01110011011100000111011101110101",
		"01100111011100010111010101110110",
		"01110111011100100110101001101000",
		"01100001011010100110110101110000",
		"01101010100000000101101001110011",
		"10000001011111100111110101111111",
		"01110101011101110110010101111001",
		"01110100011011110111000101110101",
		"01101111011000000110011001111001",
		"01101101011100100110111101100001",
		"01011000011111000110100110000000",
		"01111111011100000110111001111000",
		"01110001011101101000000010000100",
		"01110010011101100110001001011100",
		"01111000011011010111001001110011",
		"01101111011000100110010101110110",
		"01101010011100010110011101101000",
		"10000100011111000111110001111001",
		"01111101011101101000011001101010",
		"01011111011100010110111001101100",
		"01111001011011110110011001010010",
		"01111000011101100111011001111001",
		"01110101011001010101100001101101",
		"01110011011100110111000001110100",
		"10010010100010000111101101110001",
		"01101110011110011000000110001101",
		"01100010011011010111001101101011",
		"01111000011100010110011101100101",
		"01110100011101100111100101110010",
		"01101000010110010101101001100111",
		"10001101011110110111001001111000",
		"10101000100100111001001001111001",
		"01110111011100111000100010010001",
		"01100001011001110111011101101010",
		"01111001011101110110110101100011",
		"01110100011101110111011001110110",
		"01101010010110100110101101110000",
		"01110101011101110111001101110010",
		"10101011101010001001110101111010",
		"01110101011111100111001110010000",
		"01101100011010010111000101110110",
		"01110010011101100111001101100110",
		"01111000011100010111100001110001",
		"01111100011110000111010001110101",
		"01101111011100100111110101110101",
		"10011110101011011001100010000111",
		"01101110011101101000000110001010",
		"01110110011101110111011101110101",
		"01110111011101010111010101110000",
		"01110101011110000111011001111000",
		"01110111011101100111100101111100",
		"01100111010110110111100110001000",
		"10010101101000101001010110001011",
		"01101000011011101010000010000111",
		"01110000011011110111010101101111",
		"01110110011101010111001001101100",
		"01111001011100110111000101111001",
		"01101010011100110111010001110111",
		"01100101010110110111000010000001",
		"10010010101000111001000110001000",
		"01011111011000110110111110000101",
		"01101111011011110110111001101100",
		"01110101011110010110111101110010",
		"01110010011110010111100001110010",
		"01110010011010100110110101110111",
		"01111000011010000110111010000101",
		"10000101101011001001010010010010",
		"01010110010111100110011010100011",
		"01101111011011100111000001011111",
		"01110011011101110111011101110001",
		"01110101011110100111100001110101",
		"01101011011001100111000101111000",
		"01111010011101101000010101110101",
		"01110000101010011001001001110110",
		"01011101010111010101011101111010",
		"01101011011010100111001101101001",
		"01110110011101100111000001111001",
		"01110000011101010111000001111001",
		"01101011010111100110011101110001",
		"01110011100010110111010101110110",
		"10000010100101101001000110001001",
		"01101110011010110101101001100110",
		"01110111011111010111010001110100",
		"01111001011100100111000001111010",
		"01111000011101100111010001110101",
		"01101000010100010101110101110100",
		"01110101011110001000010010000101",
		"01100011100100011000110010000100",
		"01110100011110000111000101011000",
		"01111001011110001000001110001110",
		"01110011011101100111101010000001",
		"01110100011101010111010001110100",
		"10001000011011000101001001101001",
		"01111001100001111001000101111011",
		"10000000011101011000011001111000",
		"10010110011111100110100110011001",
		"01111111011110000111010110001000",
		"01110100011110010111110110001010",
		"01110111011101110111100001110100",
		"10001100011110000101001101110000",
		"10001100100100001000101110010111",
		"01101110011110000111010110000011",
		"10011100101011001010011110011000",
		"01110101011110101000110110010010",
		"01111001011110110111110010000000",
		"01111111011100100111010001110101",
		"10011011101000001010001110000001",
		"01111111100100001000010010001010",
		"10001010100010010111110110000000",
		"10001101101001010110111001110101",
		"01101110011001111001011010100010",
		"01111001011110010111100110001000",
		"01111010011101010111001001110100",
		"10001000101001101100011010000101",
		"01011111011101001000010110000110",
		"01111010011101110101001000111111",
		"10011000101001101001010101111011",
		"01110000011001011000010110011111",
		"01110010011101110111011001111011",
		"01101010011101110111101001110111",
		"10000010100011011000110001101100",
		"10000011011110001000010001111111",
		"10000101011010001000001110010010",
		"10000110011100101001100101111110",
		"01101011011011100110011001111010",
		"01110111011110110111010001110101",
		"01110000011100110111001001110010",
		"01110101011100110111010001101110",
		"01100110011100010111100001101001",
		"01110000011101000110011001101100",
		"01111101011111010111100001010111",
		"01110000011010110111010001110010",
		"01110101011100100111100101110011",
		"01110010011110000111100001110110",
		"01101000011010110110011101110001",
		"01011001010011010110101101101000",
		"01100001011010000110110001101000",
		"01101011011001100110000101011000",
		"01111001011101000111100101101110",
		"01110100011110010111011101111001",
		"01110110011101000111100001110011",
		"01110011011101100111001101110110",
		"01101011011010110110111101101111",
		"01110001011010010110100101101101",
		"01101111011100000111001101101110",
		"01110011011101000111001101110000",
		"01110100011101100111011101110110",
		"01110001011100010111010001110110",
		"01110111011101100111001001110110",
		"01111001011100010111100001110101",
		"01111010011101110111000001110100",
		"01110100011100000111000101110001",
		"01110100011101110111011101110011",
		"01110011011100010111010001110011",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"10000011000000000000000000000000",
		"01110110011100100111001001110111",
		"01111001011110000111100101111010",
		"01110100011100010111010101110100",
		"01111001011100100111001001111000",
		"01111010011101110111001101110110",
		"01111000011110000111101001110010",
		"01111010011101010111000101111001",
		"01110100011100100111011101111001",
		"01110111011101100111100001110111",
		"01110111011011110111011101110011",
		"01111110011101100111001001101111",
		"01111000011100110111001110000010",
		"01110100011110000111001101110010",
		"01110001011100110111010001110111",
		"01110010011101110111001001110101",
		"01110011011100110111011001110100",
		"10000011011111111000001101110100",
		"10001010011101110111101010000110",
		"01101111011100101000000001111101",
		"01110000011101000111010001110010",
		"01111001011100100111100101111010",
		"01110110011100100111000101110010",
		"01111101011100100111100001111001",
		"10010111100101011001110010000000",
		"10000111100100001010001110001111",
		"01110100011100111000100110010110",
		"01101101011011100110111101101110",
		"01110101011110000111001101110010",
		"01110110011101100111010101110111",
		"10000110100011110111010001101111",
		"10100110100110001001101010000110",
		"10010101101110001001000010101000",
		"01111101100100101001101110100000",
		"01011111011000000110110001110111",
		"01110111011100010111011001100110",
		"01110111011101110111100101110100",
		"01111111011110000111110001110011",
		"10011100011111100111101010001100",
		"01111110100000001000100010001111",
		"10000011100000101000010110011010",
		"01101100011101100111111110001101",
		"01110011011101110111001101100011",
		"01110111011100100111001101110110",
		"10001000011111010111101110000010",
		"01110001100110011001010101110111",
		"10000000011101100111110101111100",
		"01110100011111010111010010000100",
		"01011111011011100111001001110000",
		"01110011011100010111001101100000",
		"01111001011111000111011001110111",
		"01110010100100011000100010011001",
		"10000110011011100111010110011100",
		"01101110011110111001101101101110",
		"01101100011111010110010001111110",
		"01011001100111011000000001101100",
		"01110101011100010111001001011110",
		"01111001011100110111010101110100",
		"10000111011110011000000110010111",
		"10000000100110110110111010000011",
		"01111000011101100111000001101110",
		"10100001011001111000011101110011",
		"10000001011111010111001110001001",
		"01110101011100100110011101011011",
		"01111000011101100111000001110100",
		"01110010011001011001111110001001",
		"01101100100010011001010001110010",
		"10010110100011110111011001111010",
		"01110110100011000111101110001110",
		"01111110100010110111010101111011",
		"01110110011100010110100101011010",
		"01111011011011110111011101111001",
		"01111110101100111001101101101101",
		"10000000011101010110111101111110",
		"01101000011100100110110001111101",
		"01110011100000001001101101111011",
		"01110100011101001000000110000110",
		"01111000011110100111000101011010",
		"01110010011101110111010101110111",
		"01110101100000001000000001101111",
		"01100011010111010110101001101100",
		"01101000011001000101110101100001",
		"10011100011100110110001101110011",
		"01110100011111101000101101110100",
		"01110100011110000111110101101110",
		"01100110011101100111001101111001",
		"01011010010101000110010001100101",
		"01100011011010000110100101101010",
		"01100110011001100110100001101000",
		"10010101011001010110101001110010",
		"01100111011110111000111101111110",
		"01110111100011101010001010000101",
		"01100101011110010111011101110011",
		"01011100010011010100001101000101",
		"10010010011011010110101101101101",
		"01101001011111001010001001111010",
		"01101111011010010111011101110110",
		"01111001100000011000111001101111",
		"10001001101010001011000110111001",
		"01101000011101010111100001110011",
		"10000100011010000101010001010111",
		"10001101100000100110111101110000",
		"01110111100000011001000001111100",
		"01110100100011010110101101111110",
		"10001101011100110110111110001111",
		"01111001100110001001110010010000",
		"01110111011100010111011001110101",
		"01111100101000011010000010001001",
		"10001000011111011000000110001100",
		"10000101011111101000011101111000",
		"10000000011011110110101001111100",
		"01101001011001110110111101101100",
		"10000000100110111010011010100101",
		"10011001011100110111001001111000",
		"01111111100111101000010010011101",
		"10001011100000001001111001101110",
		"01110011100011101010000110010110",
		"10001010011101001100011101111101",
		"10001111101000001011101101101101",
		"01111101101011111100000010100000",
		"10010011100000000111001101110100",
		"10010010100101001000101010010011",
		"10001100101100011000110101111111",
		"10010010011110011000110110001101",
		"01111011011111100110011001110101",
		"01110000011111110111010101111011",
		"01111101100100111100100110001101",
		"10000000011101110111001001110001",
		"10101100100101111010111110010101",
		"10000000100100110111100101111111",
		"01101111100001011000001010110110",
		"10001110011110011001101110000000",
		"10100001100100101000100101110100",
		"01110111011110101010100010101111",
		"01101100011100100111011101110100",
		"10001100011110001000101010001111",
		"10000000101000001001101010001011",
		"10001010011111011010011101111100",
		"01101100100010011000111110001100",
		"10001111100111111000110110000010",
		"01111010100001001010100110000100",
		"10000001100000000111001001110111",
		"10111100100111101001011110010010",
		"10101100100010101001110110010111",
		"10000101011011100111101010000110",
		"10011000100001100110110101111010",
		"10001000100011111001110110100000",
		"01110100011110011000011110010100",
		"10000010100000110111100001110101",
		"10000101100010111000000110000011",
		"10000111100000011001100001100110",
		"01101100011111111000101001110001",
		"10111100100011011010010010000111",
		"10011111100100111000110001111101",
		"01110101011101111000011010000111",
		"10000010011111110111011101110110",
		"10100011100111111000010110001110",
		"01111111100000001001101110100011",
		"01110010011110000111101001111011",
		"01111000100011010111000101111110",
		"10000011100011001000000010010100",
		"01110011011100011000000010000110",
		"01110110011110010111000101110010",
		"10010011011111110111011001111001",
		"10010010011011111001011101111001",
		"01101110011100100110101010001101",
		"10101011101001010110111110001001",
		"10010001100111001001111110010001",
		"01110110011101010111111110001100",
		"01101010011100100111010101110111",
		"01101111011001110110000101101101",
		"01110111011111111000101101111001",
		"01101011111111110110010010100000",
		"10000100101001101010101001110010",
		"10000000100000001000111010000000",
		"01110011011110001000100110010111",
		"01101111011101000111011101110100",
		"01101010011011110110111001110001",
		"01101000011001110101110001011110",
		"10010101100010110111010101110100",
		"01100101011011100111111110001000",
		"01110010011001010110010101100100",
		"01111000011111000111011001111000",
		"01111000011110000111001101110111",
		"01110000011110010111000001110110",
		"01110001011101000111011101101110",
		"01101100011011100110111001110000",
		"01110010011011010110110001101110",
		"01110101011100110111001101110100",
		"01111000011100010111010101110001",
		"01110001011101010111010001110100",
		"01110100011110000111100101111000",
		"01111010011100010111011101110110",
		"01110110011101000111100101111000",
		"01110111011101100111010001110010",
		"01110110011101100111011001110110",
		"01110101011100010111100001110110",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"01010011000000000000000000000000",
		"01110101011101000111000101110100",
		"01110110011100100111001001110000",
		"01111001011101100111011001110001",
		"01111001011100110111100101110111",
		"01110111011101010111001001110100",
		"01110110011100110111100001110011",
		"01111000011100110111011001111001",
		"01110110011110100111100001111001",
		"01110110011110010111001001110011",
		"01110010011110010111001001110011",
		"01111001011100100111001101110010",
		"01110011011101110111000101110100",
		"01110111011101010111001001110001",
		"01110111011110000111100101110011",
		"01110001011100110111100001111000",
		"01110100011101100111100001110001",
		"01110111011100010111010101110100",
		"01101101011100100111010101111101",
		"01110001011011110111000001110000",
		"01110101011101010111000101111000",
		"01110111011100100111010101110010",
		"01110001011110010111001001110010",
		"10000001100000101000010001110111",
		"10011110100100001000000110001100",
		"10011000101100111000110010101000",
		"10010010100100111001100110011001",
		"01110000011010100111000110011101",
		"01110100011101000111011101110111",
		"01110111011100010111010101111000",
		"10001011100010111000110101111001",
		"10101001101001011000111110010100",
		"10011111100110101010100010101100",
		"10010001101010101000100010111111",
		"01100100011101000111010101110110",
		"01110001011101100111001001101111",
		"01111101011110010111100101110101",
		"10001110100101011001101010010000",
		"10010001100010101000011101111111",
		"10000110011111001000100010010000",
		"10011111011111000111001110100011",
		"01101111011101100111010101110110",
		"01110010011110000111010001101110",
		"10000100011101010111010001110001",
		"01111001100010011000001010000001",
		"10000111100101111001011110000010",
		"10000101011101101010000101110111",
		"01101000101001010111000110001100",
		"01111001011110111000110110000101",
		"01110010011101110111010101110011",
		"10000000011101010111101001110011",
		"10001010100010011001101010001010",
		"01110101011101111000011010010010",
		"10000111100101100111000110001010",
		"10001000011010101000101101111000",
		"01110011011011100110100001111111",
		"01110001011101010110111101110000",
		"01111011011100110111010001110110",
		"01111001011101010111111110010101",
		"01111001100011110110110101110001",
		"01111010100000101000000110000101",
		"10000100100111110111111010001000",
		"01100010101010001000001101111110",
		"01110001011100010110111101011110",
		"10000101011101010111011101110010",
		"10011000100100011000101110101001",
		"01100100011100111000001010001100",
		"10100010100110010110100101101010",
		"10001111011111111000100010010110",
		"01101100101011111000000010101001",
		"01110010011100100111000101011000",
		"10010100011101010111000001110111",
		"01110010100000010111000010001010",
		"01100111011001100110011001101101",
		"01110101011101111000100001100010",
		"10001001100011101000100110010001",
		"10000001100110110111010010001011",
		"01110000011100110111001001100100",
		"10011000011100100111000001110010",
		"01101110011101100110111110001111",
		"01110100011001110110101001110001",
		"10010011100100111001011110000100",
		"01111010011111101001100001110110",
		"01110010100100100111000011000011",
		"01110110011100000111100001100001",
		"10000000011100000111000101110111",
		"01111000011100010111000101110110",
		"01111000101000000111001101101111",
		"10000110100111110111111010010100",
		"01110111100001110111011010001110",
		"01100101011010000110100101111010",
		"01110001011100010111100001101100",
		"01110111011110010111010001110100",
		"01110110011101000110111101101000",
		"01111011011100100111001001110011",
		"01110000100100001001111010001100",
		"01111100100010110111101110001010",
		"01100111010101010110100101110001",
		"01110010011110010111101101110000",
		"01111100011110010111011001110110",
		"01101111011010110110011001101011",
		"01110011011110110111101001110100",
		"10000001100001011000010010010101",
		"01101000100000100111111001111100",
		"01110010011010010111111001101111",
		"01110100011100010110111101110110",
		"01111000011101010111100101110001",
		"01101110011110000111000001111001",
		"10000000011100100110111101101000",
		"10001100100001110111001010000110",
		"01111100011011100111111001111111",
		"10100010100100101001000010100111",
		"01110110011100100110111010010000",
		"01111111011111110111010001111000",
		"01101111011100101001000010010101",
		"01111111011110110111101001100111",
		"01110100011101001011111101110001",
		"10010010100110000111110001100110",
		"10100111100101101000000010001100",
		"01110011011100100110100110100111",
		"10010010011110100111100101110100",
		"10001010011101011000010110100001",
		"01101001011010000110011101110001",
		"01100101011001000110011001100111",
		"10100000011101101001100101110110",
		"10011110100001010111111001110010",
		"01110011011011110110010101101110",
		"10100100011110010111001101110010",
		"01111000101010001001100010001110",
		"01101111011011010110100101111010",
		"10001001011001110110101101101000",
		"10000000011111111000001010100000",
		"01111111101001101001111101111110",
		"01110011011101110110110001100110",
		"10010111011011010111000001111001",
		"01110101011101111010000010001101",
		"01110000100000110111010110000001",
		"01110101011110010111110001110011",
		"10001111100010101001011101111110",
		"10011000011110011000110001110010",
		"01110110011100110110110101110010",
		"10010110011100100111001101111001",
		"10010011101011101001100010011001",
		"01111001011111111010110110001111",
		"01110101100001100111001101100011",
		"01111011100110111000101001111110",
		"10001110100000011001001110111110",
		"01110001011101000110111101110010",
		"10001110011110000111011101110100",
		"10011001100100010111000010001101",
		"01110101011101100110011110001011",
		"01111101011100010111010101110101",
		"10101100100011110111101110000111",
		"01110010100000100111000101101101",
		"01110000011100100111011001100110",
		"10001011011111110111010101111000",
		"10001101100011000111100110000110",
		"10001010011101111000001101111101",
		"10001000011011100110111101101111",
		"01111111011101011001010001111110",
		"01110000100001110111010110011000",
		"01111010011101000110111101101101",
		"10010100100000010111011001110011",
		"10010101100011111000110010011010",
		"10010110100010111000101110000000",
		"01111000011011011001000101101000",
		"01111111101110010111001001101000",
		"01101101011011100111010010000100",
		"01111000011101010111001001101111",
		"10001010011110010111100101110001",
		"10011110101000101000010010011000",
		"10011111100111100111111110001011",
		"01111101101100011001110010000000",
		"01110011011011011010000010100101",
		"01110011011110001000000101111100",
		"01110010011100010111001001110000",
		"01101011011110100111010001111001",
		"10100110100110011000000101111000",
		"10101100101111001100000111001011",
		"10100011100011111100100111010011",
		"10100010100111001001110110101101",
		"01110001011101110111001001111010",
		"01110111011100010111011101110101",
		"01111000011100010111011101111000",
		"01110111011110010111011001110000",
		"10001010011111100111010001111000",
		"01111110100001001000110101111100",
		"01111011100001101000100110010000",
		"01111001011110010111001101111001",
		"01111010011100010111000101110101",
		"01111000011101100111100101111001",
		"01110010011110000111100101110101",
		"01110101011101000111001001110111",
		"01111000011100100111000101110111",
		"01110110011100100111010101110011",
		"01110100011101010111101001110100",
		"01110001011110010111001001110110",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"10001001000000000000000000000000",
		"01111001011101000111001001110011",
		"01110110011110010111100101111000",
		"01110111011110010111001101110011",
		"01111000011101010111000101111000",
		"01111000011100010111010101110001",
		"01110100011101000111100001111001",
		"01110001011101010111011101111010",
		"01110001011101100111100101110100",
		"01100111011011100111010101110110",
		"01101001011100100111001101101100",
		"01100011011101010110110101100011",
		"01110101011100100110111101101000",
		"01110101011100000111000101110011",
		"01111001011100100111011101111001",
		"01110110011110010111010001110010",
		"01100110011100000111100001110110",
		"01011110010111100110101101100110",
		"01100101011010100110001101011000",
		"01101111011010100110111001100100",
		"01101111011011100110111001101100",
		"01110001011100010111100101111000",
		"01110100011100110111001101110011",
		"01101011011011110111011101110011",
		"01011000010110100101010001010111",
		"01100000010110010011111001001110",
		"01110010011001100110100101100001",
		"01110110011101010111001101110111",
		"01110001011101100111100101110001",
		"01111001011100100111010101110111",
		"01110001011001100111011101111000",
		"01101111011000110110011001100010",
		"01110100011101010111110101110100",
		"10010011011101111000000010000010",
		"10010010100111111001111110011101",
		"01111001011100100111011010001110",
		"01111001011110000111001001110011",
		"01110100011100000111110001111110",
		"10000111011110111000001001111000",
		"01111101011111010110100110010000",
		"10001011100010010111111110001011",
		"10011001100010100111110110000011",
		"01110100011011100111001101111101",
		"01101110011100100111100001111000",
		"01111100011111001000110001111101",
		"01110010011100101000100001111101",
		"01100000011001110110100001101111",
		"01110100011010000110111001100111",
		"10011101100000000111001101110100",
		"01111001011110100111000101111101",
		"01110011011100100111000001110010",
		"10000110100001001001000110000010",
		"01110100011011101000001101111110",
		"01100111011000100110100001100011",
		"01111101011100110111011101100101",
		"10011011100011101000010001111111",
		"01110110011110110111101110001100",
		"01110101011111000111010101110010",
		"10001010100001111001000001111001",
		"01111111011011111000100001110001",
		"01101010011001010110100001101011",
		"01110000100000000111001001100111",
		"10001011011010001000100101110110",
		"01110110011100001000111010001101",
		"01101100011101100111011001110010",
		"01111010011110000111111001101000",
		"01111011011011100111010101111111",
		"01101010010111010110111101101110",
		"01111011100011010111100110001001",
		"10000111011111101000100010000111",
		"01110001011100100111000001101101",
		"01101001011011110111001001111000",
		"01111001011011010110011101101000",
		"01111100011100111000100101111001",
		"01101111010100010110010110010001",
		"10010001011111110111111101100110",
		"01100011100001101000101101110111",
		"01110100011011110110011001101010",
		"01101111011011000110111101111001",
		"10001110100011111000000001100100",
		"01111011101101001010101110010001",
		"10100101010101100100110010110110",
		"01111101100000001000111110100011",
		"01011100011101000110111001110110",
		"01110101011100100110001101010101",
		"01100011011001100111001101111000",
		"10110000100100101000000101011111",
		"10011101101001110111110010101011",
		"10000110011001110111011011011101",
		"10001000011110110111100010001111",
		"01101111100011101010100110001100",
		"01110100011010110110110001110110",
		"01101000011011100111010101110110",
		"10011010100111101000100101110101",
		"10100100101000011001110010001100",
		"10100100011101100110110010101101",
		"01111111100011001000101010001101",
		"01110100100101001010010010011011",
		"01101111011101000111000101100100",
		"01101111011011000111011001111000",
		"10011000100100111010001010011111",
		"10010011100010011000011110000110",
		"10000111100000010110101110101111",
		"10100101100000001010001010010100",
		"01110011100011001000010010000110",
		"01111000011010000111001001101000",
		"01111110011110100111100101110100",
		"10010011100100101000010010001111",
		"10100001100011111001100010010000",
		"10001001100001000110011110001000",
		"10010001011111111010000110100001",
		"01111011100110100111010101110000",
		"01110000011100110110010101001000",
		"01101001011100010111011101110110",
		"10010111100000100111000101011010",
		"01111100011111111000011110010111",
		"10100011100011110111111010001010",
		"10000011100000111001001110001111",
		"01111010011110011000111110011100",
		"01110100011010000110100101100101",
		"01011100011101000111100101111001",
		"10001111011110100111010001101011",
		"01111110100001111000111010010010",
		"10001100101001000111111101110111",
		"01101011100110001000111110001111",
		"01110011011101001001000101111100",
		"01101111011011100101111101100001",
		"01101100011110000111001001110110",
		"10001000100001000111110101111010",
		"01110101011011001000110110001010",
		"10000000100001101001100010100010",
		"01110111011100010110101010010010",
		"01101110011000101000011110000011",
		"01110010011101010101110101100010",
		"01111110011100000111011001110010",
		"01111000100011101000100101110101",
		"01110111011010110110101001101100",
		"01110101100100000110101101011110",
		"01110001011101010110111001110110",
		"01011101010110011000000001101111",
		"01110010011100110110100001100101",
		"01111100011110000111010101110110",
		"01101010011100100110100001111001",
		"01110101011010100111000101101001",
		"01110111011100010110010001101111",
		"01110001011111101000101110001111",
		"01100001011010110111101001110011",
		"01111000011101100110100101100101",
		"01101111011101110111000101110001",
		"01101000011001000111010001101110",
		"01110110011100110111100110001101",
		"01111011011011010110011101110000",
		"10000010011101101000010001100111",
		"01110111011110110111111010000111",
		"01110111011110000110101101101101",
		"01110010011110100111100101111000",
		"01101101011010100110011101101101",
		"01101111011011110110110101110010",
		"01101011011011000111000001101000",
		"10011101011101110111111001101110",
		"01110001100000111001010001111001",
		"01110010011110000110111101101111",
		"01110001011110010111011101110010",
		"01111100011111000110101001110100",
		"01110001011101101000001110000011",
		"01110001011110110111000101101110",
		"10001011100100110111101010001100",
		"01100111011010101000100110001000",
		"01111000011110010111010101101111",
		"01110100011110000111011001110010",
		"01111011011110010111001101110000",
		"10110111011100111000101101111000",
		"01110010100000110111011101110000",
		"10000011011110010111010010001000",
		"01110011011110000111101101111000",
		"01110110011101010111100101110011",
		"01110111011101000111100101110111",
		"01100111011010110111001101111000",
		"01110111100001100111000101100101",
		"10000110100000101000001001110001",
		"01100010011100100111001001110011",
		"01110001011100000110010101101010",
		"01110011011101000111000001110001",
		"01110001011101000111010001110011",
		"01100111011100000111010101111010",
		"01011110010111100101110101100100",
		"01010111010011100101100101100011",
		"01011010010101000101100101011001",
		"01110101011010100110011001100110",
		"01111000011110000111000101110110",
		"01110100011101000111011101110100",
		"01110010011011110111100001111000",
		"01110010011100010111011001101111",
		"01101111011001100111011001101110",
		"01110101011011110111001001110011",
		"01110101011100000110110101110101",
		"01110101011100010111001001110111",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"11111110000000000000000000000000",
		"01110101011100010111000001110010",
		"01110101011100010111100101110111",
		"01110010011101000111001101110010",
		"01110100011101000111011101110010",
		"01110101011101110111010001110010",
		"01110011011101000111001001110100",
		"01110111011100100111011101111000",
		"01110100011101110111011101110111",
		"01110001011101100111001001111001",
		"01110010011100010111100001110001",
		"01110110011101100111010001110010",
		"01110001011100100111100001111001",
		"01111000011110000111100001110011",
		"01111010011101100111001001110001",
		"01110100011100110111000101111001",
		"01110110011100110111010101111010",
		"01101011011011000111001101110111",
		"01110000011010110110101001101101",
		"01110111011111100111111001110101",
		"01110010011100010110110001101110",
		"01110011011101010111011001101111",
		"01110110011101110111011101110001",
		"01110010011101100110101101110101",
		"01101101011100000111010001101111",
		"10001111011110100111110101111011",
		"10001000100110001000101001110100",
		"01110001100001011001100010010011",
		"01111001011110100111110001111110",
		"01110010011100100111100001110111",
		"01101110011001010110000101101101",
		"10101001011101010110111101100111",
		"11010111011110000111000110100111",
		"10001011101111101001001010000000",
		"10001110100000011001011101101011",
		"01110011011110001000101110011100",
		"01101111011101000111011001111001",
		"01110100011000100110001001011111",
		"10001000100111110111011001110011",
		"01101100011101011000001001111111",
		"01110100100001011001000110000011",
		"10001100100011100111101010100100",
		"01110010011111011001001010010100",
		"01100110011110010111100101111000",
		"01110111011101010111001001100000",
		"01111000011101100111011001111001",
		"01111000100010110111100010000101",
		"10011010100000010111110101110111",
		"10001011100011110111000110001001",
		"01110110100001001001011110100101",
		"01101000011101010111100101110110",
		"01111001011111000110110001001110",
		"01111101100101100111010010110001",
		"01100100100001110110101010000010",
		"01110101100000110111110110000011",
		"10010111100101011000100001111110",
		"01111000011111101010110010101011",
		"01100101011110000111000101110111",
		"01101101011110100110101001000010",
		"10000000100000111000100101111110",
		"01110000011100110111001101111000",
		"10001100011110011000000001111110",
		"10110001011100111000100010010111",
		"01110101100010001011001111000110",
		"01100010011100000111001001110011",
		"01110100100000010110111001010100",
		"10010001011111100110110001111100",
		"01100110011100000111001001111111",
		"01110101100000110111100101100111",
		"10011000100111111011011001110101",
		"01110111100010111011101111010111",
		"01100111011101000111011101111000",
		"10010100011011100111001001110000",
		"10000110100101011010000110011100",
		"01110100011110101000011010011000",
		"01101111011010100110100001101101",
		"10111110011010010111001001110000",
		"01111010100101011110000011110011",
		"01100010011101000111100101111010",
		"10010000100101100111011001110100",
		"10001011100001001000100110010010",
		"01110010100001101010111010001011",
		"01101001011100100110111101110100",
		"01110011010111000110100001100111",
		"01110001100010111101001011000101",
		"01101100011101110111011101110100",
		"10001110101001010111010101110111",
		"10001110101000010111110110000100",
		"10001000011101001001011110001111",
		"01100111011010010110010001101100",
		"00111110010101000101111101101111",
		"01110101100011000111010100101011",
		"01110010011101000111010101110001",
		"10100001011100101001011110000100",
		"10010110100000010111111101111010",
		"01101011011101111001101010101000",
		"10000011011100110111001001100101",
		"01011001011011010110111110000111",
		"01110011011100110101111100111000",
		"01110101011101010111001001110111",
		"10000001011101010111001110000000",
		"10000001100110011000000010000000",
		"01110111011111010111111010001010",
		"01100111011010010110100101110000",
		"01110100100010100111000101111100",
		"01110100011100100101100101110111",
		"01101111011100110111100101111000",
		"01101111011110110110111101110011",
		"10000010100001111000111001111001",
		"01101101011011100111110010001110",
		"01111001100111010111000101111010",
		"10001101011001011000100101110111",
		"01101110011011010110011010010010",
		"01110100011100110111011101110101",
		"01101000011011110111001001101111",
		"01110110100000000110100001110000",
		"01111010011011110111101101111011",
		"10000000011001100111100101101000",
		"10001111101001010111100110011001",
		"01110000011010110110101101111101",
		"01111010011010110111001001111001",
		"01101101101001111000100101111101",
		"01110001011101010111011101110100",
		"01111000011010010110100001100111",
		"01111111100110101001000101111111",
		"10001100011100001000010001111111",
		"01110101011100000110010001111010",
		"01111011011101110111100001111001",
		"10010010101101101001000110100111",
		"01111110011110110111010101110101",
		"01111111011111110111100101110011",
		"10000001011010011000100101111111",
		"10010000100011000111011101110001",
		"01110110011011110110100110001110",
		"01111100011111100111010101110110",
		"01110110100110100111010010100101",
		"10000110100011100111010010101000",
		"01111101011011101000100110000000",
		"01110011100010000111001001110000",
		"10010101100000101001001010011100",
		"01110100011100010111000110001001",
		"10000010100000000111010101111000",
		"01111000100100011010011101111111",
		"10001010100000001010000110010110",
		"01110101011100111000100001111000",
		"10010110100010011000111110001011",
		"10000111101011000111110001111111",
		"01111001011100111000000001111100",
		"01111001011100000111001101110100",
		"10100100100100100111101110010000",
		"10001011011111101000010010001001",
		"01111110100000100111101001111100",
		"01111110100000001000110001110010",
		"10000111100110111001101010011110",
		"01110100011101000111110010000100",
		"01111010011100100111100001111001",
		"10000011011100010110110110010100",
		"01111110011100010111111101111011",
		"01111110100010001000000010000000",
		"10001101100110100111011110000111",
		"10010010100010110111101110000101",
		"01110110011101001000000010001011",
		"01111111011110000111011101111000",
		"01101101100001111001000010000111",
		"10000001101001000111011110011001",
		"01110010100000110111001010000110",
		"01110111011011110111011110001011",
		"10000101100000000111100110001101",
		"01110011011101000111100010000000",
		"01111001011101010111011001110100",
		"01111011011111000111110101111011",
		"10001011100001111010011110001010",
		"10100001101000011010011110001101",
		"10000001101000101010110110000000",
		"01111111100010110111011010001001",
		"01110100011110100111000101111010",
		"01111001011110010111011001110101",
		"01111001011111010111010110000001",
		"10101011100111101001111001111000",
		"10111000011111111011000110101010",
		"10001100100101011010000110101111",
		"10001011100011011000111010000001",
		"01110001011101000111011110000001",
		"01110111011110010111011101110101",
		"01100111011011010111011001110110",
		"10000001011101010110100001100101",
		"10001011011111010111111110001100",
		"01110010011010010111000001111011",
		"01110111011100110111011101111010",
		"01110101011101010111001001110111",
		"01110110011110010111001101110111",
		"01110110011101000111010001110001",
		"01110010011101100111000101110010",
		"01110010011100110111000101111001",
		"01110100011101010111011101110010",
		"01110011011101100111011101110100",
		"01110010011100010111010101110010",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"01101111000000000000000000000000",
		"01110011011101000111001001110101",
		"01110010011100100111011001110101",
		"01110101011100010111000001110110",
		"01110011011100110111001001111001",
		"01110100011110010111010101110110",
		"01111001011110010111000101110110",
		"01110111011101010111001001110100",
		"01110001011110010111001101111000",
		"01111111011111010111100001111001",
		"01111011011110100111110010000000",
		"01111000011110001000001010000111",
		"01111110011111000111011101110101",
		"01111100011110100111101001111000",
		"01110111011100100111001001111001",
		"01110111011100000111000001111001",
		"10001100011111100111001001111010",
		"10010100100100111000100110001111",
		"10000011100010111000101010010011",
		"10001100100001001000010110000011",
		"01111110100001101000111110000111",
		"01110111011110000111000101110110",
		"01111000011100110111010001110010",
		"10000111100000010111010001110110",
		"10010000100011111001000110001000",
		"10001100100011001001000010001100",
		"10001101100010000111110110000011",
		"10001101100001100111111101111001",
		"01110011011101010110110010000001",
		"01110100011110010111001001110111",
		"01110101011111010111100001111011",
		"01111101100001110111000110000001",
		"10000010100001011000001101111111",
		"10000000100000011001000110010011",
		"10001011100011001000011110000101",
		"01111010011110000110101101100000",
		"01101111011100100111010101110110",
		"01101100011100100110100001110110",
		"01101011100011110111101110000110",
		"01101101100000010110110001110101",
		"10011010100011011000010001110011",
		"10011110011100101000101010000110",
		"01111010011101110111001001111111",
		"01101111011110000111010001111000",
		"01110101011000110110110001110101",
		"01101110011010000111010101110111",
		"01110110011010000110011101110000",
		"01101000011001100110111101101010",
		"10001000011100100111010101101111",
		"01110110011110110111010110001110",
		"01101111011110000111000101111001",
		"01111111011000100111011001110011",
		"01111010011100000111010101110011",
		"01110001011100110110001101110001",
		"01101000011010000110101101100111",
		"01110101011011100111010001101001",
		"01110101011100110111000010001000",
		"01101101011101010111010101110101",
		"01110000011011100111010001110111",
		"01101111011100000111100001110010",
		"01011100011000000111010001101001",
		"01100000010110100110110001101000",
		"01100101011011010111000101101010",
		"01101111011011000110010101100001",
		"01110100011100110111101001111001",
		"01111100011011100110100110000010",
		"01110000011001010110101101110000",
		"01100111011011110101110001101100",
		"01100100010110100101100101011101",
		"01101101011011010111101001101110",
		"01110000011001010101101101101000",
		"01101011011100110111001101110100",
		"01111111011100010110110001110010",
		"01101110011101110110111110000000",
		"01011100011001110111010001101101",
		"01101000011001010110011101100100",
		"01110100011001000111000101110010",
		"01110011011001100101100001110001",
		"01110010011100100111100101110100",
		"10010110011101000111110001110101",
		"01110111100000101001101110000110",
		"01011100011101001001011110010001",
		"01111010011001110110011101110101",
		"10011011011011101000010101111001",
		"01110100010110000101001001111000",
		"01101011011101100111011101110000",
		"10100010100011010111110001110011",
		"10100001100001111000111010010011",
		"01101010011011111001001010010001",
		"01100011011011010111010001111100",
		"10111101101001011001001001111001",
		"01110001010110000110000110011001",
		"01101111011101010111000101110010",
		"10001001101010011000100101110001",
		"01111001100011110111100101110110",
		"10000100011011111001011010010000",
		"10000100011100100110110001111101",
		"10110101100011101001011101111010",
		"01110010010110100101100110011001",
		"01110010011100010111011101110101",
		"01111010100100101000101001011110",
		"10100100100101101000111110001101",
		"01111111011100110111100110001011",
		"01111101011110000110010110001101",
		"10010001100011111000101001111001",
		"01110001011001100111111010010000",
		"01110001011110100111001001111000",
		"10010000100100000111000001011001",
		"10010001100010010111111110010001",
		"01111011100101111000101110010101",
		"01111010011110101000001001111011",
		"10000001011110111000110110000110",
		"01110111011000111000110010000110",
		"01101000011101010111011101110100",
		"10010110101001011000010101011011",
		"10110100100100011001110010001110",
		"01111101100010000111100001111001",
		"10001010100010100111001010000001",
		"01111000100001001000100101111011",
		"01101111011000111000100010000001",
		"01110000011101110111100001111000",
		"10001000100001011000001101011000",
		"10101100101011011001111110010110",
		"01110111100100001000100110000101",
		"10000110100000001000100001110101",
		"10000111100010111000010110000011",
		"01110101011010111000101010000110",
		"01110011011101100111001001110010",
		"10011110100000000111001001100000",
		"01111101100011111001000110001001",
		"01111001011101001001101010110000",
		"01111001100011001000101110001111",
		"10001001011101110111110101111010",
		"01110101011100101000001110000100",
		"01110010011110100111010101110110",
		"10001001100100010111100101110011",
		"10101010101000011001110001111000",
		"10001011100110011000011110100011",
		"10000101100001001000101110000011",
		"10001101100111001000100001111111",
		"01110011011100100110100001110011",
		"01110011011101010111100001110111",
		"10011101011101010111010001101110",
		"10010100101001101001111101101110",
		"10001110101000110111111110011111",
		"01111100100101001000001110001000",
		"10000000011110001001000110011010",
		"01110110011101000110110101101101",
		"01110101011100100111010101110101",
		"01111100011010100110011001101000",
		"10001100100011001000101110100111",
		"10001001100110111001010110100101",
		"10001111101000111001111110001000",
		"01101110100000110111001010010111",
		"01110111011101010110111001110000",
		"01110101011100110111100001110110",
		"01110101010111100110011101101011",
		"01101010100111101000011001111111",
		"10100111011010011001001010010001",
		"01111111011110110111011010000101",
		"01100100011010011000011110001100",
		"01111001011101100111100001100110",
		"01111000011101110111011101110000",
		"01100111011010110111001101110001",
		"01101111011010010111000001101010",
		"01110101011110110111010001110110",
		"10010010100101010111011101110100",
		"01101101011011100111011010000001",
		"01110001011110010111001001101101",
		"01110001011101000111100001110111",
		"01110010011101000111001101111001",
		"01011000011000000110010001101010",
		"01101111011010000110001101100101",
		"01101101011101010111100101111011",
		"01110010011100100111000101110000",
		"01110101011100100111100001110010",
		"01110110011100100111010101110010",
		"01110010011101110111000101110110",
		"01110101011100100111001101110101",
		"01101010011100000110110101110111",
		"01101111011100110111001101101111",
		"01110011011101010111100101110011",
		"01111000011100010111011001110000",
		"01111001011110010111010101110011",
		"01110010011101100111001101110010",
		"01111000011100010111010001110010",
		"01110011011101110111001101110010",
		"01110001011101100111100001111001",
		"01110001011101000111001001111001",
		"01110010011110000111000001110001",
		"01110110011100100111000101110010",
		"01110100011101110111100001111001",
		"01110111011101110111000101110101",
		"01111000011101000111010001111000",
		"01110011011101100111001101110011",
		"01110010011100100111010001110100",
		"01110111011110010111000101110011",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"11010100000000000000000000000000",
		"01111001011101000111001101111001",
		"01110101011110010111000101110100",
		"01110100011100110111001001110001",
		"01110111011110000111011101110101",
		"01110000011101110111001001110001",
		"01110110011101000111000101110010",
		"01110011011110010111001001110110",
		"01111001011101110111100101110011",
		"01110001011101100111000101111001",
		"01110111011101110111101001111001",
		"01110100011110000111000101110100",
		"01110100011110010111011001110110",
		"01110001011100110111000101110111",
		"01110001011110010111100001110001",
		"01110101011101010111000101111000",
		"01110101011101110111010001111000",
		"01110100011100000111000001110111",
		"01110100011100010111010001110101",
		"01110010011101100111001001110101",
		"01110000011110010111001001110001",
		"01110011011101100111001101110101",
		"01110100011100010111001101111001",
		"01110101011101110111101001111000",
		"01101001011010000111001101110010",
		"01101101011011110110100101101011",
		"01110100011101110110111001110001",
		"01110111011110000111011001110111",
		"01110111011100110111100101110111",
		"01110001011100100111001101110101",
		"01101011011011000111010001110110",
		"01011100010101110101111101101001",
		"01100101011001010110100001100100",
		"01101010011010110110011101100110",
		"01110100011100010111010101101111",
		"01110101011101100111011101110001",
		"01110100011101000111100101110010",
		"10000100011110100111110001110010",
		"01110111011101101001010110010010",
		"01110001011100101000000110001011",
		"01100101011011100110111001110011",
		"01101111011010010110011101011011",
		"01110111011110000111000101110000",
		"10000110011101000111010001110101",
		"10010000100101011000110101111111",
		"10101110100011101000111010011010",
		"01111100011110110111010010010010",
		"01111001011111111000101010000101",
		"01100101011101001000011101110011",
		"01111000011110000111000101101101",
		"10010011011111110111010101111001",
		"10011001100011000111110110001010",
		"01111011100011101000110101111011",
		"10001001011011011000110110001111",
		"01110111101000111000101010001011",
		"10000000100000111000110110100100",
		"01110100011110010111001001111000",
		"10010101100000000111101001110010",
		"10100101100011101000101110001100",
		"10010010011111111001000110011000",
		"10011000100010100110111110011100",
		"10000010100111101000001010001000",
		"10001100100100100111010110010101",
		"01110101011101100110101001110010",
		"10001111100000000111110101110111",
		"10000110100100111000101010010001",
		"10000010011110001000110010000111",
		"10010100101010010111100110100011",
		"10010100100101111011010110001111",
		"10000011100100011001011101110110",
		"10000000011101010111100001111100",
		"10010001100010110111111101110010",
		"10000110100011101000110110001111",
		"01100110011101101001000101111000",
		"10001100100010001001100001100111",
		"10100001100010111000011010110100",
		"01110111100111001001101010101011",
		"01110010011110110111011101101011",
		"10010001100110110111110001110101",
		"10010001100001100111111010001101",
		"10010100101101101001000001101110",
		"10100110101100111000100010000110",
		"10000010101010011000111110001011",
		"01110000100111001001001010101010",
		"01110111011100110110111001100101",
		"10100000100110010111111001110101",
		"10101001011110011000100010011110",
		"10011000011100010111000011011010",
		"10101011011011010101000001011101",
		"01111010101000001001011110100111",
		"01101110101010111000111001111001",
		"01110011011111010111011001100101",
		"10011000100010100111011001111000",
		"10000000101100101000001110001110",
		"01110000100001100111000001101000",
		"01111010011100010101100101001111",
		"01100111011100110111101010001110",
		"01101100011110011010000010010000",
		"01110011011101010111110001111010",
		"10001001100000000111101001110100",
		"01110110011101101001000110001001",
		"01100011011101000111000101111010",
		"01110001011100010110001001011001",
		"11000011100011011000100110001001",
		"10010100100010100111000110011111",
		"01110010011110000110111001110010",
		"10000011011101110111000001110110",
		"01110001011110100111001101110000",
		"01100111011100010110101101101100",
		"10001100011001100110110001011100",
		"01111011101000111100000001011111",
		"10010111101000011000111110010110",
		"01110010011011100110000001101011",
		"01101101011101110111001101110100",
		"10100111011101110110111001111101",
		"01011010011010000111000001111001",
		"10001011010110010111110101101110",
		"10010010011110111001100001111000",
		"01110010011100101001010110011000",
		"01110001011011110110011101101000",
		"01101010011100010111011001110001",
		"01101111011101011000000010000010",
		"01101101011001110111001001110100",
		"10001000100001011000000110000110",
		"01101110100011010111011001110111",
		"01110110100000000111010110001100",
		"01110000011101110111110110000010",
		"01101110011101110111010001110001",
		"01101100011001110111111101111101",
		"01111000011101000110111101101110",
		"01110001011100101000001101101110",
		"01110100011101100111011101110010",
		"01011101011101011000000001110011",
		"01111001011101010111011101101101",
		"01101101011111000111011001110110",
		"01100111011011000110111101110100",
		"01110001011000000111001101110011",
		"01101000011111100110111001110100",
		"01110010011001000110101001101000",
		"01010101010110100110111001110001",
		"01110111011110010111010101101111",
		"01100110011100010111010001110001",
		"01100110010110110110001001011110",
		"01101110011011100110111001110011",
		"01100110011110110111010001111011",
		"01100111010110100110000101100000",
		"01100010010100010101111001011010",
		"01110100011101010110110001101110",
		"01101000011100000111010101110100",
		"01011101010111010110001101011010",
		"01101111011101010110111101110100",
		"01101000010111110110010001110001",
		"01100110011010000110100101110100",
		"01010111010100000101101001100101",
		"01110110011100110111000001110100",
		"01100010011010010111010101111010",
		"10000001011100010111000101011110",
		"01100111011101010111001001110111",
		"01110000011101110110000001111101",
		"01110101011010110110101001110111",
		"01011001010100010101011101100011",
		"01110001011100110111010101101111",
		"01100011011100110111011001111001",
		"10011100100011110111101001110010",
		"01100111011011100110111001011101",
		"01111010011011100110001001100100",
		"01101000011011010111001001110000",
		"01010110010101000101000101011001",
		"01110001011100010111010001101111",
		"01110111011101010111001101110101",
		"10001110100101111001101101111111",
		"01111101100000010111010110001011",
		"01111001011110111000111101110000",
		"01101101011010001000010101110011",
		"01011011011001010110100001101011",
		"01110100011101100110111101101110",
		"01110111011101010111010001110111",
		"10000100011100110111011010000100",
		"10110110100101111010000110010100",
		"10011010101000001001100010101110",
		"01111111100100011001000010011000",
		"01110001011101010111010101110000",
		"01110001011110000111011101110001",
		"01111001011110000111100101110110",
		"01111011011000100110100001101111",
		"10000101100011011000110010000100",
		"10011101100101011001010110000001",
		"10010110100101101001011110001100",
		"01110100100000100111100001110110",
		"01110001011110010111011001110000",
		"01110111011110100111011001110011",
		"01110011011101110111000101110010",
		"01111001011111000111010101111000",
		"01111100100000011000011001111011",
		"10000011100001001000000101111111",
		"01110100100000001000000001111011",
		"01111001011100110111001101110110",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"01111000011101100111000101110001",
		"01110011011101000111001001111001",
		"01110110011100000111001001110100",
		"01110111011101000111011101110101",
		"01110001011101010111100101111000",
		"01110010011101000111011001111010",
		"01110001011100100111001001110011",
		"01111001011100100111011101111000",
		"01111010011100100111100101110001",
		"01110010011101000111100101111000",
		"01110110011101110111100001110011",
		"01111000011100010111010101110110",
		"01110100011100010111011101110011",
		"01110011011101110111010001111001",
		"01110110011100100111010101110010",
		"01110011011110010111000101110110",
		"01110000011100000111100001110100",
		"01110000011100110111000101110000",
		"01110011011101010110111001101110",
		"01110101011100110111001001110101",
		"01110011011101000111001001111001",
		"01110010011101010111100101110110",
		"01110001011100100111001001110001",
		"01110100011110010111010101111000",
		"01110110011101010111100101110011",
		"01110001100011101000001101110110",
		"10000010100010000111110101110010",
		"01111000011100010111010001110101",
		"01110110011100100111010101110100",
		"01110010011011000111000101110011",
		"10001011100111001001000010000101",
		"10100001110001010110010011011101",
		"01110010101110011000101110110011",
		"01111110100100001000000110100111",
		"01111000011111001000010110000110",
		"01110000011101100111100001110110",
		"10000010011011000110101101110101",
		"10100011011011011000011001110001",
		"01111111100010011000000010010000",
		"10001000011011011010000010000111",
		"01101101011101110111111010010111",
		"01111000011101101000111010000011",
		"01110110011100100111011001110100",
		"01110011011011110110111001101111",
		"01110101011110101000001001111010",
		"10001111100000001000000010011011",
		"10011111011011111000110101111110",
		"10011101011101010111011110000001",
		"01110010011101111001001101110001",
		"01110000011100010111011101110001",
		"01101100011011100111010101110010",
		"01101101100001000111001110100111",
		"10001110011000000111110101101110",
		"01110111100010000110111001111011",
		"10101000011111001001010001110010",
		"01110011011101100111111010011001",
		"01111100011100110111010001110001",
		"10011011100101101000100101111001",
		"01111001100010101000101101110001",
		"01110011011011101000101110000110",
		"10010010100010110111011110001111",
		"10001010100001011000111110000010",
		"01111111100010011001000110110011",
		"01110010011101100111010001110110",
		"01111110100100110111011101110110",
		"10000111011110001000101110010000",
		"01100101011101110111110001101001",
		"10000001011101101000101101111100",
		"10011010100010011000111010000001",
		"01110010100100001001011110011100",
		"01101110011100110111011001110100",
		"01110101100001000111010010010010",
		"10000011100110001000100101111010",
		"01011110011101010111100110011011",
		"10011101100100110111011001101100",
		"10010011100100001001001110010000",
		"01110101011110100111001001110110",
		"01110001011100010111011001110101",
		"11000110100010101000111010000001",
		"10001011100100101010001010100110",
		"01111110101101001001101010001111",
		"01110101011010010111000001111001",
		"10010110100100010111100110000000",
		"01110101100001100111100110010111",
		"01111110011110010111011101110100",
		"10100100011100001010010001111000",
		"10000111011111001000110001101101",
		"10000111100001101001111010001101",
		"10011100011100111000011101111101",
		"10110001101000011011000110001001",
		"01110000011101110111100110111100",
		"01111011011101110111100101110000",
		"01111011100110001000001001110010",
		"10010000011011101000000001111110",
		"10011001011101111010100010011001",
		"01110110011111010110111110001000",
		"10011100100010000110101010101100",
		"01111000011101010111110110010000",
		"01110111011101000111011101110000",
		"01101101011110010111100001100101",
		"10011100100000010110100101101011",
		"10000011100010101001100110001110",
		"01111101011101001000001110000010",
		"01100011011001110111010001101011",
		"01110011011101010111101101100111",
		"01110011011101100111010101111001",
		"01110101011100110110011101101001",
		"01111001011101011000011001110001",
		"10000001100110101001000010001101",
		"01111001100001000111011101111001",
		"01101010011101000111001101110000",
		"01110110011100000111101001100101",
		"01111010011101010111001001110110",
		"01110100011101010110101101101000",
		"10000101100100100111110101110101",
		"01111110100001101000101010011001",
		"01100111011100111000100010001000",
		"10000100011011000111000101101101",
		"01110100011011110110100001101010",
		"01110101011101100111010101110011",
		"10110011011100000111000101110010",
		"10001100100000111001110110001011",
		"01110000100000111000100110010001",
		"01110111011001100111011110000110",
		"10001110011101010111101101110101",
		"01111000011100000110001010000111",
		"01101100011101000111010101110011",
		"01110100100110000111010001101100",
		"10010111100101101001001101111111",
		"01110110011101011000010110001101",
		"01110001011101100110110101110011",
		"10010000011100110110111110000011",
		"01111001011101000110001001110001",
		"01100111011101000111001101110010",
		"01101111100001101010010001101110",
		"01110011100011101000111010000011",
		"01110010011100100111001110000011",
		"10000000100010001000001101111110",
		"10100110101000100110101101110100",
		"01110110011100100110010001101011",
		"01100110011100010111001101111000",
		"10101001011110010111011001101111",
		"01110101100100100111110010001000",
		"10000010011001011000001001111110",
		"10001010011110000111100101101010",
		"10001010100011001011000110011101",
		"01110111011101100110100101100111",
		"01101010011101100111011001110101",
		"10100011101000000111010001110110",
		"01111101011010111001010101110110",
		"01110011011101111000001001101000",
		"01111111011111101001000101110010",
		"01110110100011110110111110001110",
		"01110100011101100110111101100010",
		"01110101011100010111001101110001",
		"10001010100011010111100001111101",
		"10000011011110100111100001101110",
		"01111111100001010111100101111101",
		"01110100011111110111110001110100",
		"01111101011110111000101001101011",
		"01110111011100100111000001101110",
		"01110100011110010111011001111001",
		"01101011011010000110101101110100",
		"10000010011111000111111010011111",
		"10000101011110111001011110000101",
		"10010101101000010111101010000110",
		"10000100100000001000000110001000",
		"01110101011101010111001001101110",
		"01101011011101100111011101110110",
		"01110000011001100101110001100110",
		"10100011011111011000001110011111",
		"10001010101010001001001010010101",
		"10111111100111100110011111001000",
		"01110001011100000111001010001000",
		"01110001011100100111010101101100",
		"01111001011100110111100101110011",
		"01110001011100000110001001101101",
		"10101011101001000111000101110000",
		"10100110101001100111110010001101",
		"10001001100001011010101110100000",
		"01101101011100110110111101111011",
		"01110100011101100111100101110100",
		"01110110011101110111100001110011",
		"01110101011010110111010101110111",
		"01110011011011000111000101110100",
		"01100111011010110111010001110100",
		"01101111011100010111000101101010",
		"01110001011101000111000001101010",
		"01110110011101100111010001110110",
		"01110010011110000111101001110011",
		"01111010011101110111010001110011",
		"01111001011101010111100001110100",
		"01110001011101100111100101110101",
		"01110101011110010111001101110101",
		"01110011011101100111000101110011",
		"01111001011110010111100001110111",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"01100011000000000000000000000000",
		"01110010011110010111010101110110",
		"01110101011101000111011101110100",
		"01110010011100100111011101110110",
		"01111001011100110111100101110001",
		"01111001011110100111100001110011",
		"01110100011100100111010101110111",
		"01110101011101110111000101110100",
		"01110100011100010111001001110010",
		"01110010011101010111100001110110",
		"01110001011100110111010101110011",
		"01110101011110000111100001110010",
		"01110100011101010111100001110000",
		"01110101011101010111011101110010",
		"01110101011110010111011001110111",
		"01111001011110000111100001111000",
		"01110011011100100111100001111001",
		"01110100011100010111001001110101",
		"01110011011101010111000101110101",
		"01110101011101010111001001110010",
		"01110001011101000111001001110100",
		"01110111011101110111011001110100",
		"01110100011101110111011101110111",
		"01110010011110010111000101111001",
		"01101101011100100111001101110001",
		"01100110011010100110011101101010",
		"01110001011101000110111101101000",
		"01110001011101010111000101110010",
		"01110111011110010111011101110110",
		"01110100011100110111100101110100",
		"01110011011110000111010001110100",
		"01101110011011000110110001101110",
		"01110110011101000111000101101111",
		"01100100011011100110111101101111",
		"01110011011010110110011101101000",
		"01110111011101010111001101110010",
		"01110100011100110111010001110110",
		"01101011011100000111010001111001",
		"10111100011010010110111001101101",
		"10001001011001111000111010001111",
		"01110101011100100111001001101010",
		"01101001011001110111000001110100",
		"01110110011101010111001001101101",
		"01110101011100110111001001111001",
		"01101111011001110101111001101100",
		"10011010011100001001010101110100",
		"10001001100011111001101101111110",
		"01110111101000101001000110010111",
		"01101110011100010111011010010111",
		"01110101011100000111000001101101",
		"01101101011100100111000001110111",
		"01101111011100000101101001100100",
		"01111010011110100111100001110100",
		"10011011100011111001100110010011",
		"10000001100001101000101110011011",
		"01111100011101010111010110001111",
		"01110100011011010111000101101111",
		"01100100011100000111011101110111",
		"01100111011110010110111101100001",
		"01110111011110010111100010101000",
		"10000011100100001000010101100101",
		"01111111100011000111111010001110",
		"01111011011101111010110001101101",
		"01110011011100010110111101111001",
		"01100111011010100111001101110011",
		"01110101101001000111011101100110",
		"10000001100011100111111001111100",
		"10011011100010100111110001111111",
		"10000010100011011000101001111110",
		"01110100100001100110110010001000",
		"01110111011100110110111001110100",
		"01101000011011010110111101111000",
		"01110111101000000111011001101110",
		"01111101100000101000010110001000",
		"01101101011101110110011010000010",
		"10001110100001010111011001111110",
		"01110100011111010111100110000010",
		"01111000011101010111001001100111",
		"01100011011000000110110101110101",
		"10010111100001010111111101101110",
		"10010110101000011001011010110010",
		"10011101100001001001010110011100",
		"01111110100100001001110010010001",
		"01110010101001011001110010111011",
		"01110001011100110110100101100111",
		"01100110011010000111000001111000",
		"10011100101011011001100110001110",
		"10010111100100111001011110010111",
		"10010111100011001000010001110101",
		"10010101100101011000110010001110",
		"10100110101001101010101010001000",
		"01110111011011110110101001100000",
		"01101110011001110111001001111001",
		"10100000011111111001001010110011",
		"10000101100001000111100010001111",
		"10010001100010011000111101111001",
		"10011110100010001000101010011110",
		"01101010100001111001110010011000",
		"01110110011011000110000001010011",
		"01110100011100000111011001110100",
		"10000010101000010111111110010010",
		"10000000100000110111110101110101",
		"10001010011111001000111010000001",
		"01111111100001101001010010001111",
		"01011110011111101001010010010001",
		"01110111011100010110100101010001",
		"01110100011011000111100101111000",
		"10000010100001000111111010000011",
		"10001001100000110111101010001000",
		"10001101011011100111101101110100",
		"10001100100000001001110110001100",
		"01100110011110110111000110000100",
		"01110100011011100110110001010100",
		"01110000011100000111001101110010",
		"01111100011101001000001110000001",
		"10001011100001110111000110001111",
		"01111010011111000111001101110111",
		"01101011100000111000111110001011",
		"01100001100001000111000101111001",
		"01111010011100110110010001010110",
		"01101010011100100111100101110101",
		"10001011011100000111000001100100",
		"01110000100011000111100110010001",
		"10010000011101111000010010000111",
		"01110001011111101000000101111011",
		"01100001011011110111010001110100",
		"01110101011101100110110101011001",
		"01101000011101000111011101110100",
		"01111101100010010110011101100011",
		"10010100101010010111000001110001",
		"01111110100011010110101001101000",
		"01101111011100100111111101111011",
		"01011011011011010111010010000011",
		"01110011011100010110110101010110",
		"01101000011101000111001001110101",
		"10001010011111010110100101100011",
		"01101000011011100110111001111001",
		"01100100011010000110110001110101",
		"10000010011101000110011101110101",
		"01100111011010010111000001111110",
		"01110011011101000110110101101101",
		"01100101011100100111000101110001",
		"01101111011101010111111101101101",
		"01011011011001110110110001110010",
		"01100100011011000110101101011001",
		"01111001011100010111100001110111",
		"01110100011011110110100001110000",
		"01111001011101110111101010000100",
		"01101110011101110111000101110001",
		"01110100011111100111100001101110",
		"01100011011011010111000101110001",
		"01100100010111000101111001100011",
		"01110100011010110110100001110000",
		"01110101011010000111011101110100",
		"01110101011100110111010010000100",
		"01110110011101100111101001111001",
		"01110100011100100110011001101110",
		"01110110100001110110111110001011",
		"01011101011110010110100001111001",
		"01101000011011110110111001101100",
		"10000101011100100110110101111000",
		"01110110011101100111011110000000",
		"01110001011101000111000001110010",
		"01101111011011000110100101100111",
		"01110000011100100110100010000001",
		"01101101011111110111000101101111",
		"01111110011110000111001001110011",
		"10000110100111001000101001111100",
		"01110100011100010111010010000101",
		"01110001011110010111011101110010",
		"10000011011111000111100101110111",
		"10000000100010110110101110010001",
		"10000001011001110111000101110010",
		"10001001100010001000101010000110",
		"10001011100011111000011110001111",
		"01110010011100100111000001101011",
		"01110001011100010111011001111000",
		"10010000100100001001110001110111",
		"10100000101001011001001010011101",
		"10010011101010101001100110100101",
		"10001101100100101001010110011101",
		"01111011011101101001001010011100",
		"01110011011101000111011001101110",
		"01110111011100110111001001110110",
		"10100001100110101000111001111110",
		"10100001101001011010110010100010",
		"10010111101110001010010010101111",
		"10001101101001001001011010011100",
		"01111010011101111000100010001101",
		"01111001011101010111010001110111",
		"01110011011110100111100001110110",
		"01111001011101100111001101111000",
		"01110011011101110111011101111000",
		"01111011011101100110100101111010",
		"01110000011101000111001001110001",
		"01111000011101100111100001111000",
		"00000000000000000000000000000000"
    );

    signal rom_index: std_logic_vector (11 downto 0);
begin
    rom_index <= (in_rom_neuron_index & in_rom_input_index); -- combine the neuron and input index to adress the array
    out_data_rom <= rom_arr(to_integer(unsigned(rom_index)));
end RTL;
