library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
    port (
        clk, reset:             in std_logic;
        in_rom_input_index:     in std_logic_vector(7 downto 0); -- the given rom input index
        in_rom_neuron_index:    in std_logic_vector(3 downto 0); -- the given neuron index
        out_weights:            out std_logic_vector(31 downto 0) -- the output datastream
    );
end ROM;

architecture RTL of ROM is 
    type t_rom_arr is array (0 to 2500) of std_logic_vector (31 downto 0);
    constant rom_arr: t_rom_arr := (
        -- here follows the generated array allocation
        2500 => "01110001011101010111100001111010",
        2499 => "01110101011011010111011001110101",
        2498 => "01111001011110000111011001110101",
        2497 => "01110011011100010111100101110001",
        2496 => "01110100011100100111011101110011",
        2495 => "01110100011110010111010001111001",
        2494 => "01110111011101010111100101110001",
        2493 => "01110111011101000111100101111001",
        2492 => "01110111011100010110110001101110",
        2491 => "01110000011100010110110001101110",
        2490 => "01101110011011100110101101110110",
        2489 => "01110100011011100111000001101111",
        2488 => "01110101011101100111011001110001",
        2487 => "01110110011100010111011101110100",
        2486 => "01110001011110000111100001111000",
        2485 => "01110111011011010110011001100110",
        2484 => "01100101010110110101101101100100",
        2483 => "01011011010110110110000101011110",
        2482 => "01100010010111010110011101100110",
        2481 => "01101010011011000110111101110000",
        2480 => "01110111011101000111011101111001",
        2479 => "01110101011101100111001101110001",
        2478 => "01110100011010000110010101011011",
        2477 => "01100000011101001000001110000011",
        2476 => "10001101100110001001101110011110",
        2475 => "01110101100011001000011101111011",
        2474 => "01101100011011100111001001110010",
        2473 => "01110101011101000111100001110101",
        2472 => "01110001011100100111010001101101",
        2471 => "01101110011101000110100101100110",
        2470 => "01101110011100001000111001110010",
        2469 => "01111110100010011000011110000101",
        2468 => "10011001100110011000111110000101",
        2467 => "10001101011110000110100001100000",
        2466 => "01110011011110010111011001110011",
        2465 => "01110100011100010110111101101000",
        2464 => "01110111100001000111011001111001",
        2463 => "10000101011100111000101101111110",
        2462 => "10000001011110011010100110000010",
        2461 => "01110111100010101000100110001100",
        2460 => "01111111100011001000000001011110",
        2459 => "01110110011101010111011101110111",
        2458 => "01110100011111010111001001101000",
        2457 => "01101110011111110111101101111001",
        2456 => "01110010011100110110111001111100",
        2455 => "01111011011100000111010010010011",
        2454 => "10001101100010100111110101111000",
        2453 => "10010011100011001000011001110101",
        2452 => "01110110011100010111011001110110",
        2451 => "01110101011101000111001001101110",
        2450 => "01101101100101011000100001111111",
        2449 => "10000000011111101000000101101101",
        2448 => "10000000011100101000100010100111",
        2447 => "10010011100101111001001110010100",
        2446 => "10001010100100001001010010000011",
        2445 => "01101111011110010111010101110110",
        2444 => "01111001011100110111000101110111",
        2443 => "01111110100110011000110110000001",
        2442 => "01101110100000110111111101101001",
        2441 => "01101101011011000110100010011010",
        2440 => "10011100100011010111101110010010",
        2439 => "10010010100100111000001101111110",
        2438 => "01101101011100010111011001110010",
        2437 => "01110011011110000111000001111011",
        2436 => "10000011100100100111010101101111",
        2435 => "01110001011101010111101001110101",
        2434 => "01110000011010000110000001101110",
        2433 => "01111010101001111001011110011001",
        2432 => "10000101100011000111111110000001",
        2431 => "01110000011101010111100101111000",
        2430 => "01110101011100010110111101111101",
        2429 => "10000011100010110111100110001101",
        2428 => "10000000011101001001110101110010",
        2427 => "01101000011000100101111001110100",
        2426 => "10000010101100001001011101111001",
        2425 => "10001111100110011001000110000101",
        2424 => "01110101011101000111100101110010",
        2423 => "01110010011101000110101110000010",
        2422 => "10001000100011001000100110010001",
        2421 => "10000000100000101000001001101011",
        2420 => "01101010010111000101100001101011",
        2419 => "10010111100011001001000110011001",
        2418 => "10001111100100001001010010001000",
        2417 => "01110010011100110111100001110100",
        2416 => "01110110011100000111110010011001",
        2415 => "10010010100010001000001110010001",
        2414 => "01110011011111100111000001100010",
        2413 => "01011010010011100110010001110011",
        2412 => "01101100100111111001000010010010",
        2411 => "10011101011101001001100110001010",
        2410 => "01100111011100000111100101110110",
        2409 => "01111001011101111000010010100000",
        2408 => "10011000100000111000111010000111",
        2407 => "01110100011110000111000101011001",
        2406 => "01011001010110000110110110101111",
        2405 => "10011110011011101000111010000110",
        2404 => "10100001100010001001001001110000",
        2403 => "01101010011100100111011101110110",
        2402 => "01110110011100011000000110011011",
        2401 => "10010111100011010111110101101001",
        2400 => "01111001011110010110111001011011",
        2399 => "01010011010110010110011010000010",
        2398 => "01111010100111010111111110001001",
        2397 => "10010110100111010111100110000100",
        2396 => "01110101011100110111101001110001",
        2395 => "01111000011011100111000110101110",
        2394 => "10010011100101001001000110010000",
        2393 => "10001101011101000111001101011110",
        2392 => "01011001011000011000011010101000",
        2391 => "10000100100000110111111001111111",
        2390 => "10001110101000010111011101110000",
        2389 => "01110100011101000111010001111001",
        2388 => "01110100011001110110011110010010",
        2387 => "10001101100101001010000110001111",
        2386 => "10000010011010010111001101011100",
        2385 => "01011011011011001000001001101000",
        2384 => "10001000011111110111001010001111",
        2383 => "10010000100001110110111001101101",
        2382 => "01110101011101100111001101111000",
        2381 => "01110110011001010110000110100000",
        2380 => "10011000100101001000100110001110",
        2379 => "01110011100101101011011001111111",
        2378 => "01101110100011111000110101111001",
        2377 => "10001101011100111001001001111001",
        2376 => "01111100011110011000011101110011",
        2375 => "01111001011101110111000101110010",
        2374 => "01110010011001110101111110100011",
        2373 => "10011011011100110111011110001110",
        2372 => "10011001100100111001000010001000",
        2371 => "01100010011101011001111101110010",
        2370 => "01110010100100100111110101110000",
        2369 => "01110101011100010111011101110001",
        2368 => "01111110011100100111100101110011",
        2367 => "01110111011001100101011010001111",
        2366 => "10101000100011001001000010010000",
        2365 => "01110111100001111000111110101100",
        2364 => "10001101100011100110111010001100",
        2363 => "01110100011110101000111110000001",
        2362 => "01111010011110100111010101101100",
        2361 => "01110111011100010111010101111001",
        2360 => "01110001011001000101110101110001",
        2359 => "10010001011100110111110001111000",
        2358 => "10001000100100101001010101110000",
        2357 => "01110011011111001000011001110100",
        2356 => "10001000100000101000100001110000",
        2355 => "10000111100000110111011101110001",
        2354 => "01110100011110000111001001110011",
        2353 => "01110110011011000101110001011110",
        2352 => "01110011100111111001100110001000",
        2351 => "01111101100011101000000010001101",
        2350 => "01110010100011111001000001101111",
        2349 => "01110111011111000110100001111111",
        2348 => "01111110100000010111000001101111",
        2347 => "01111000011101110111001101110110",
        2346 => "01110010011100000110011101100110",
        2345 => "01101100011110101000000001110010",
        2344 => "10001001100101011001001110000101",
        2343 => "10000001100100001001000101110100",
        2342 => "10010011100110011000010010000001",
        2341 => "01111011011101010110010101110101",
        2340 => "01110101011101100111011101110111",
        2339 => "01111001011101000111000101101100",
        2338 => "01110101011110100111010001111001",
        2337 => "10000001100010111001011110000111",
        2336 => "10011000100001011001011010001001",
        2335 => "10100000011111111000011001111000",
        2334 => "01110110011001110110101001110010",
        2333 => "01110111011100010111100001110001",
        2332 => "01110001011101000111011101110100",
        2331 => "01110011011011010110100101110010",
        2330 => "01110010011101101000101010001111",
        2329 => "10000011100100011000111101111010",
        2328 => "01111100011110110111010001110101",
        2327 => "01100111011011010110111001111001",
        2326 => "01111000011100100111011101110010",
        2325 => "01110001011101010111010101111001",
        2324 => "01110011011100100111000101101110",
        2323 => "01110001011100000110110101101100",
        2322 => "01100111011010110110111001110110",
        2321 => "01110011011100100111010101110101",
        2320 => "01110101011100010111100001111000",
        2319 => "01111001011101010111100001110010",
        2318 => "01110010011110010111010001110101",
        2317 => "01110001011100010111011101110111",
        2316 => "01111000011110010111101001111100",
        2315 => "01110100011100000111100001111001",
        2314 => "01110101011100010111011101111001",
        2313 => "01110110011101100111001101110010",
        2312 => "01111000011101110111010101110110",
        2311 => "01110101011101100111100101110010",
        2310 => "01111001011100010111010101110111",
        2309 => "01110001011110010111100001110110",
        2308 => "01110101011100110111011001110101",
        2307 => "01110100011110000111001101110010",
        2306 => "01111000011101010111011001110001",
        2305 => "01110110011101000111001001111000",
        2304 => "01010000000000000000000000000000",
        2244 => "01110011011100010111010001110011",
        2243 => "01110100011101110111011101110011",
        2242 => "01110100011100000111000101110001",
        2241 => "01111010011101110111000001110100",
        2240 => "01111001011100010111100001110101",
        2239 => "01110111011101100111001001110110",
        2238 => "01110001011100010111010001110110",
        2237 => "01110100011101100111011101110110",
        2236 => "01110011011101000111001101110000",
        2235 => "01101111011100000111001101101110",
        2234 => "01110001011010010110100101101101",
        2233 => "01101011011010110110111101101111",
        2232 => "01110011011101100111001101110110",
        2231 => "01110110011101000111100001110011",
        2230 => "01110100011110010111011101111001",
        2229 => "01111001011101000111100101101110",
        2228 => "01101011011001100110000101011000",
        2227 => "01100001011010000110110001101000",
        2226 => "01011001010011010110101101101000",
        2225 => "01101000011010110110011101110001",
        2224 => "01110010011110000111100001110110",
        2223 => "01110101011100100111100101110011",
        2222 => "01110000011010110111010001110010",
        2221 => "01111101011111010111100001010111",
        2220 => "01110000011101000110011001101100",
        2219 => "01100110011100010111100001101001",
        2218 => "01110101011100110111010001101110",
        2217 => "01110000011100110111001001110010",
        2216 => "01110111011110110111010001110101",
        2215 => "01101011011011100110011001111010",
        2214 => "10000110011100101001100101111110",
        2213 => "10000101011010001000001110010010",
        2212 => "10000011011110001000010001111111",
        2211 => "10000010100011011000110001101100",
        2210 => "01101010011101110111101001110111",
        2209 => "01110010011101110111011001111011",
        2208 => "01110000011001011000010110011111",
        2207 => "10011000101001101001010101111011",
        2206 => "01111010011101110101001000111111",
        2205 => "01011111011101001000010110000110",
        2204 => "10001000101001101100011010000101",
        2203 => "01111010011101010111001001110100",
        2202 => "01111001011110010111100110001000",
        2201 => "01101110011001111001011010100010",
        2200 => "10001101101001010110111001110101",
        2199 => "10001010100010010111110110000000",
        2198 => "01111111100100001000010010001010",
        2197 => "10011011101000001010001110000001",
        2196 => "01111111011100100111010001110101",
        2195 => "01111001011110110111110010000000",
        2194 => "01110101011110101000110110010010",
        2193 => "10011100101011001010011110011000",
        2192 => "01101110011110000111010110000011",
        2191 => "10001100100100001000101110010111",
        2190 => "10001100011110000101001101110000",
        2189 => "01110111011101110111100001110100",
        2188 => "01110100011110010111110110001010",
        2187 => "01111111011110000111010110001000",
        2186 => "10010110011111100110100110011001",
        2185 => "10000000011101011000011001111000",
        2184 => "01111001100001111001000101111011",
        2183 => "10001000011011000101001001101001",
        2182 => "01110100011101010111010001110100",
        2181 => "01110011011101100111101010000001",
        2180 => "01111001011110001000001110001110",
        2179 => "01110100011110000111000101011000",
        2178 => "01100011100100011000110010000100",
        2177 => "01110101011110001000010010000101",
        2176 => "01101000010100010101110101110100",
        2175 => "01111000011101100111010001110101",
        2174 => "01111001011100100111000001111010",
        2173 => "01110111011111010111010001110100",
        2172 => "01101110011010110101101001100110",
        2171 => "10000010100101101001000110001001",
        2170 => "01110011100010110111010101110110",
        2169 => "01101011010111100110011101110001",
        2168 => "01110000011101010111000001111001",
        2167 => "01110110011101100111000001111001",
        2166 => "01101011011010100111001101101001",
        2165 => "01011101010111010101011101111010",
        2164 => "01110000101010011001001001110110",
        2163 => "01111010011101101000010101110101",
        2162 => "01101011011001100111000101111000",
        2161 => "01110101011110100111100001110101",
        2160 => "01110011011101110111011101110001",
        2159 => "01101111011011100111000001011111",
        2158 => "01010110010111100110011010100011",
        2157 => "10000101101011001001010010010010",
        2156 => "01111000011010000110111010000101",
        2155 => "01110010011010100110110101110111",
        2154 => "01110010011110010111100001110010",
        2153 => "01110101011110010110111101110010",
        2152 => "01101111011011110110111001101100",
        2151 => "01011111011000110110111110000101",
        2150 => "10010010101000111001000110001000",
        2149 => "01100101010110110111000010000001",
        2148 => "01101010011100110111010001110111",
        2147 => "01111001011100110111000101111001",
        2146 => "01110110011101010111001001101100",
        2145 => "01110000011011110111010101101111",
        2144 => "01101000011011101010000010000111",
        2143 => "10010101101000101001010110001011",
        2142 => "01100111010110110111100110001000",
        2141 => "01110111011101100111100101111100",
        2140 => "01110101011110000111011001111000",
        2139 => "01110111011101010111010101110000",
        2138 => "01110110011101110111011101110101",
        2137 => "01101110011101101000000110001010",
        2136 => "10011110101011011001100010000111",
        2135 => "01101111011100100111110101110101",
        2134 => "01111100011110000111010001110101",
        2133 => "01111000011100010111100001110001",
        2132 => "01110010011101100111001101100110",
        2131 => "01101100011010010111000101110110",
        2130 => "01110101011111100111001110010000",
        2129 => "10101011101010001001110101111010",
        2128 => "01110101011101110111001101110010",
        2127 => "01101010010110100110101101110000",
        2126 => "01110100011101110111011001110110",
        2125 => "01111001011101110110110101100011",
        2124 => "01100001011001110111011101101010",
        2123 => "01110111011100111000100010010001",
        2122 => "10101000100100111001001001111001",
        2121 => "10001101011110110111001001111000",
        2120 => "01101000010110010101101001100111",
        2119 => "01110100011101100111100101110010",
        2118 => "01111000011100010110011101100101",
        2117 => "01100010011011010111001101101011",
        2116 => "01101110011110011000000110001101",
        2115 => "10010010100010000111101101110001",
        2114 => "01110011011100110111000001110100",
        2113 => "01110101011001010101100001101101",
        2112 => "01111000011101100111011001111001",
        2111 => "01111001011011110110011001010010",
        2110 => "01011111011100010110111001101100",
        2109 => "01111101011101101000011001101010",
        2108 => "10000100011111000111110001111001",
        2107 => "01101010011100010110011101101000",
        2106 => "01101111011000100110010101110110",
        2105 => "01111000011011010111001001110011",
        2104 => "01110010011101100110001001011100",
        2103 => "01110001011101101000000010000100",
        2102 => "01111111011100000110111001111000",
        2101 => "01011000011111000110100110000000",
        2100 => "01101101011100100110111101100001",
        2099 => "01101111011000000110011001111001",
        2098 => "01110100011011110111000101110101",
        2097 => "01110101011101110110010101111001",
        2096 => "10000001011111100111110101111111",
        2095 => "01101010100000000101101001110011",
        2094 => "01100001011010100110110101110000",
        2093 => "01110111011100100110101001101000",
        2092 => "01100111011100010111010101110110",
        2091 => "01110011011100000111011101110101",
        2090 => "01110111011011110110001101101110",
        2089 => "01111111100010101000100001111111",
        2088 => "01111101011111010110101001111100",
        2087 => "10000101011101010111101001101101",
        2086 => "01101010011100010110100001100111",
        2085 => "01111001100001001000000001111010",
        2084 => "01111010011110000111001001110111",
        2083 => "01110110011100110110100101010101",
        2082 => "01101010011011010111100101111110",
        2081 => "10000011011111001000001110001010",
        2080 => "10000111100010101001000110000011",
        2079 => "01110110011110010111001101111100",
        2078 => "01110010011111100111101001110001",
        2077 => "01110010011101110111100001110100",
        2076 => "01110011011101010111011101110000",
        2075 => "01101111011011010110101001110010",
        2074 => "01110100011001110111011010001101",
        2073 => "10000100011101000111110001110101",
        2072 => "01100010011001100110111001110000",
        2071 => "01110100011101000111100001110100",
        2070 => "01110111011100000111011001110011",
        2069 => "01111001011110000111100101110101",
        2068 => "01111001011100110111000101111000",
        2067 => "01110100011110000111011010001000",
        2066 => "10010010011111111000001101110001",
        2065 => "01110000011011010110111101110101",
        2064 => "01110100011100100111100001110100",
        2063 => "01110110011101100111100101111000",
        2062 => "01111001011100100111001101110001",
        2061 => "01110101011101000111000101111001",
        2060 => "01111010011101010111001101110100",
        2059 => "01111010011110100111011101110001",
        2058 => "01111010011110000111011001110100",
        2057 => "01110010011101110111010101111000",
        2056 => "01110111011101000111100001110011",
        2055 => "01110110011110010111010001110111",
        2054 => "01110100011100010111011101110111",
        2053 => "01111000011101110111000101110111",
        2052 => "01111000011101110111000101110001",
        2051 => "01110110011100010111000101110100",
        2050 => "01110010011110010111001001110011",
        2049 => "01111000011101000111010001110111",
        2048 => "10111001000000000000000000000000",
        1988 => "01110101011100010111100001110110",
        1987 => "01110110011101100111011001110110",
        1986 => "01110111011101100111010001110010",
        1985 => "01110110011101000111100101111000",
        1984 => "01111010011100010111011101110110",
        1983 => "01110100011110000111100101111000",
        1982 => "01110001011101010111010001110100",
        1981 => "01111000011100010111010101110001",
        1980 => "01110101011100110111001101110100",
        1979 => "01110010011011010110110001101110",
        1978 => "01101100011011100110111001110000",
        1977 => "01110001011101000111011101101110",
        1976 => "01110000011110010111000001110110",
        1975 => "01111000011110000111001101110111",
        1974 => "01111000011111000111011001111000",
        1973 => "01110010011001010110010101100100",
        1972 => "01100101011011100111111110001000",
        1971 => "10010101100010110111010101110100",
        1970 => "01101000011001110101110001011110",
        1969 => "01101010011011110110111001110001",
        1968 => "01101111011101000111011101110100",
        1967 => "01110011011110001000100110010111",
        1966 => "10000000100000001000111010000000",
        1965 => "10000100101001101010101001110010",
        1964 => "01101011111111110110010010100000",
        1963 => "01110111011111111000101101111001",
        1962 => "01101111011001110110000101101101",
        1961 => "01101010011100100111010101110111",
        1960 => "01110110011101010111111110001100",
        1959 => "10010001100111001001111110010001",
        1958 => "10101011101001010110111110001001",
        1957 => "01101110011100100110101010001101",
        1956 => "10010010011011111001011101111001",
        1955 => "10010011011111110111011001111001",
        1954 => "01110110011110010111000101110010",
        1953 => "01110011011100011000000010000110",
        1952 => "10000011100011001000000010010100",
        1951 => "01111000100011010111000101111110",
        1950 => "01110010011110000111101001111011",
        1949 => "01111111100000001001101110100011",
        1948 => "10100011100111111000010110001110",
        1947 => "10000010011111110111011101110110",
        1946 => "01110101011101111000011010000111",
        1945 => "10011111100100111000110001111101",
        1944 => "10111100100011011010010010000111",
        1943 => "01101100011111111000101001110001",
        1942 => "10000111100000011001100001100110",
        1941 => "10000101100010111000000110000011",
        1940 => "10000010100000110111100001110101",
        1939 => "01110100011110011000011110010100",
        1938 => "10001000100011111001110110100000",
        1937 => "10011000100001100110110101111010",
        1936 => "10000101011011100111101010000110",
        1935 => "10101100100010101001110110010111",
        1934 => "10111100100111101001011110010010",
        1933 => "10000001100000000111001001110111",
        1932 => "01111010100001001010100110000100",
        1931 => "10001111100111111000110110000010",
        1930 => "01101100100010011000111110001100",
        1929 => "10001010011111011010011101111100",
        1928 => "10000000101000001001101010001011",
        1927 => "10001100011110001000101010001111",
        1926 => "01101100011100100111011101110100",
        1925 => "01110111011110101010100010101111",
        1924 => "10100001100100101000100101110100",
        1923 => "10001110011110011001101110000000",
        1922 => "01101111100001011000001010110110",
        1921 => "10000000100100110111100101111111",
        1920 => "10101100100101111010111110010101",
        1919 => "10000000011101110111001001110001",
        1918 => "01111101100100111100100110001101",
        1917 => "01110000011111110111010101111011",
        1916 => "01111011011111100110011001110101",
        1915 => "10010010011110011000110110001101",
        1914 => "10001100101100011000110101111111",
        1913 => "10010010100101001000101010010011",
        1912 => "10010011100000000111001101110100",
        1911 => "01111101101011111100000010100000",
        1910 => "10001111101000001011101101101101",
        1909 => "10001010011101001100011101111101",
        1908 => "01110011100011101010000110010110",
        1907 => "10001011100000001001111001101110",
        1906 => "01111111100111101000010010011101",
        1905 => "10011001011100110111001001111000",
        1904 => "10000000100110111010011010100101",
        1903 => "01101001011001110110111101101100",
        1902 => "10000000011011110110101001111100",
        1901 => "10000101011111101000011101111000",
        1900 => "10001000011111011000000110001100",
        1899 => "01111100101000011010000010001001",
        1898 => "01110111011100010111011001110101",
        1897 => "01111001100110001001110010010000",
        1896 => "10001101011100110110111110001111",
        1895 => "01110100100011010110101101111110",
        1894 => "01110111100000011001000001111100",
        1893 => "10001101100000100110111101110000",
        1892 => "10000100011010000101010001010111",
        1891 => "01101000011101010111100001110011",
        1890 => "10001001101010001011000110111001",
        1889 => "01111001100000011000111001101111",
        1888 => "01101111011010010111011101110110",
        1887 => "01101001011111001010001001111010",
        1886 => "10010010011011010110101101101101",
        1885 => "01011100010011010100001101000101",
        1884 => "01100101011110010111011101110011",
        1883 => "01110111100011101010001010000101",
        1882 => "01100111011110111000111101111110",
        1881 => "10010101011001010110101001110010",
        1880 => "01100110011001100110100001101000",
        1879 => "01100011011010000110100101101010",
        1878 => "01011010010101000110010001100101",
        1877 => "01100110011101100111001101111001",
        1876 => "01110100011110000111110101101110",
        1875 => "01110100011111101000101101110100",
        1874 => "10011100011100110110001101110011",
        1873 => "01101000011001000101110101100001",
        1872 => "01100011010111010110101001101100",
        1871 => "01110101100000001000000001101111",
        1870 => "01110010011101110111010101110111",
        1869 => "01111000011110100111000101011010",
        1868 => "01110100011101001000000110000110",
        1867 => "01110011100000001001101101111011",
        1866 => "01101000011100100110110001111101",
        1865 => "10000000011101010110111101111110",
        1864 => "01111110101100111001101101101101",
        1863 => "01111011011011110111011101111001",
        1862 => "01110110011100010110100101011010",
        1861 => "01111110100010110111010101111011",
        1860 => "01110110100011000111101110001110",
        1859 => "10010110100011110111011001111010",
        1858 => "01101100100010011001010001110010",
        1857 => "01110010011001011001111110001001",
        1856 => "01111000011101100111000001110100",
        1855 => "01110101011100100110011101011011",
        1854 => "10000001011111010111001110001001",
        1853 => "10100001011001111000011101110011",
        1852 => "01111000011101100111000001101110",
        1851 => "10000000100110110110111010000011",
        1850 => "10000111011110011000000110010111",
        1849 => "01111001011100110111010101110100",
        1848 => "01110101011100010111001001011110",
        1847 => "01011001100111011000000001101100",
        1846 => "01101100011111010110010001111110",
        1845 => "01101110011110111001101101101110",
        1844 => "10000110011011100111010110011100",
        1843 => "01110010100100011000100010011001",
        1842 => "01111001011111000111011001110111",
        1841 => "01110011011100010111001101100000",
        1840 => "01011111011011100111001001110000",
        1839 => "01110100011111010111010010000100",
        1838 => "10000000011101100111110101111100",
        1837 => "01110001100110011001010101110111",
        1836 => "10001000011111010111101110000010",
        1835 => "01110111011100100111001101110110",
        1834 => "01110011011101110111001101100011",
        1833 => "01101100011101100111111110001101",
        1832 => "10000011100000101000010110011010",
        1831 => "01111110100000001000100010001111",
        1830 => "10011100011111100111101010001100",
        1829 => "01111111011110000111110001110011",
        1828 => "01110111011101110111100101110100",
        1827 => "01110111011100010111011001100110",
        1826 => "01011111011000000110110001110111",
        1825 => "01111101100100101001101110100000",
        1824 => "10010101101110001001000010101000",
        1823 => "10100110100110001001101010000110",
        1822 => "10000110100011110111010001101111",
        1821 => "01110110011101100111010101110111",
        1820 => "01110101011110000111001101110010",
        1819 => "01101101011011100110111101101110",
        1818 => "01110100011100111000100110010110",
        1817 => "10000111100100001010001110001111",
        1816 => "10010111100101011001110010000000",
        1815 => "01111101011100100111100001111001",
        1814 => "01110110011100100111000101110010",
        1813 => "01111001011100100111100101111010",
        1812 => "01110000011101000111010001110010",
        1811 => "01101111011100101000000001111101",
        1810 => "10001010011101110111101010000110",
        1809 => "10000011011111111000001101110100",
        1808 => "01110011011100110111011001110100",
        1807 => "01110010011101110111001001110101",
        1806 => "01110001011100110111010001110111",
        1805 => "01110100011110000111001101110010",
        1804 => "01111000011100110111001110000010",
        1803 => "01111110011101100111001001101111",
        1802 => "01110111011011110111011101110011",
        1801 => "01110111011101100111100001110111",
        1800 => "01110100011100100111011101111001",
        1799 => "01111010011101010111000101111001",
        1798 => "01111000011110000111101001110010",
        1797 => "01111010011101110111001101110110",
        1796 => "01111001011100100111001001111000",
        1795 => "01110100011100010111010101110100",
        1794 => "01111001011110000111100101111010",
        1793 => "01110110011100100111001001110111",
        1792 => "10000011000000000000000000000000",
        1732 => "01110001011110010111001001110110",
        1731 => "01110100011101010111101001110100",
        1730 => "01110110011100100111010101110011",
        1729 => "01111000011100100111000101110111",
        1728 => "01110101011101000111001001110111",
        1727 => "01110010011110000111100101110101",
        1726 => "01111000011101100111100101111001",
        1725 => "01111010011100010111000101110101",
        1724 => "01111001011110010111001101111001",
        1723 => "01111011100001101000100110010000",
        1722 => "01111110100001001000110101111100",
        1721 => "10001010011111100111010001111000",
        1720 => "01110111011110010111011001110000",
        1719 => "01111000011100010111011101111000",
        1718 => "01110111011100010111011101110101",
        1717 => "01110001011101110111001001111010",
        1716 => "10100010100111001001110110101101",
        1715 => "10100011100011111100100111010011",
        1714 => "10101100101111001100000111001011",
        1713 => "10100110100110011000000101111000",
        1712 => "01101011011110100111010001111001",
        1711 => "01110010011100010111001001110000",
        1710 => "01110011011110001000000101111100",
        1709 => "01110011011011011010000010100101",
        1708 => "01111101101100011001110010000000",
        1707 => "10011111100111100111111110001011",
        1706 => "10011110101000101000010010011000",
        1705 => "10001010011110010111100101110001",
        1704 => "01111000011101010111001001101111",
        1703 => "01101101011011100111010010000100",
        1702 => "01111111101110010111001001101000",
        1701 => "01111000011011011001000101101000",
        1700 => "10010110100010111000101110000000",
        1699 => "10010101100011111000110010011010",
        1698 => "10010100100000010111011001110011",
        1697 => "01111010011101000110111101101101",
        1696 => "01110000100001110111010110011000",
        1695 => "01111111011101011001010001111110",
        1694 => "10001000011011100110111101101111",
        1693 => "10001010011101111000001101111101",
        1692 => "10001101100011000111100110000110",
        1691 => "10001011011111110111010101111000",
        1690 => "01110000011100100111011001100110",
        1689 => "01110010100000100111000101101101",
        1688 => "10101100100011110111101110000111",
        1687 => "01111101011100010111010101110101",
        1686 => "01110101011101100110011110001011",
        1685 => "10011001100100010111000010001101",
        1684 => "10001110011110000111011101110100",
        1683 => "01110001011101000110111101110010",
        1682 => "10001110100000011001001110111110",
        1681 => "01111011100110111000101001111110",
        1680 => "01110101100001100111001101100011",
        1679 => "01111001011111111010110110001111",
        1678 => "10010011101011101001100010011001",
        1677 => "10010110011100100111001101111001",
        1676 => "01110110011100110110110101110010",
        1675 => "10011000011110011000110001110010",
        1674 => "10001111100010101001011101111110",
        1673 => "01110101011110010111110001110011",
        1672 => "01110000100000110111010110000001",
        1671 => "01110101011101111010000010001101",
        1670 => "10010111011011010111000001111001",
        1669 => "01110011011101110110110001100110",
        1668 => "01111111101001101001111101111110",
        1667 => "10000000011111111000001010100000",
        1666 => "10001001011001110110101101101000",
        1665 => "01101111011011010110100101111010",
        1664 => "01111000101010001001100010001110",
        1663 => "10100100011110010111001101110010",
        1662 => "01110011011011110110010101101110",
        1661 => "10011110100001010111111001110010",
        1660 => "10100000011101101001100101110110",
        1659 => "01100101011001000110011001100111",
        1658 => "01101001011010000110011101110001",
        1657 => "10001010011101011000010110100001",
        1656 => "10010010011110100111100101110100",
        1655 => "01110011011100100110100110100111",
        1654 => "10100111100101101000000010001100",
        1653 => "10010010100110000111110001100110",
        1652 => "01110100011101001011111101110001",
        1651 => "01111111011110110111101001100111",
        1650 => "01101111011100101001000010010101",
        1649 => "01111111011111110111010001111000",
        1648 => "01110110011100100110111010010000",
        1647 => "10100010100100101001000010100111",
        1646 => "01111100011011100111111001111111",
        1645 => "10001100100001110111001010000110",
        1644 => "10000000011100100110111101101000",
        1643 => "01101110011110000111000001111001",
        1642 => "01111000011101010111100101110001",
        1641 => "01110100011100010110111101110110",
        1640 => "01110010011010010111111001101111",
        1639 => "01101000100000100111111001111100",
        1638 => "10000001100001011000010010010101",
        1637 => "01110011011110110111101001110100",
        1636 => "01101111011010110110011001101011",
        1635 => "01111100011110010111011001110110",
        1634 => "01110010011110010111101101110000",
        1633 => "01100111010101010110100101110001",
        1632 => "01111100100010110111101110001010",
        1631 => "01110000100100001001111010001100",
        1630 => "01111011011100100111001001110011",
        1629 => "01110110011101000110111101101000",
        1628 => "01110111011110010111010001110100",
        1627 => "01110001011100010111100001101100",
        1626 => "01100101011010000110100101111010",
        1625 => "01110111100001110111011010001110",
        1624 => "10000110100111110111111010010100",
        1623 => "01111000101000000111001101101111",
        1622 => "01111000011100010111000101110110",
        1621 => "10000000011100000111000101110111",
        1620 => "01110110011100000111100001100001",
        1619 => "01110010100100100111000011000011",
        1618 => "01111010011111101001100001110110",
        1617 => "10010011100100111001011110000100",
        1616 => "01110100011001110110101001110001",
        1615 => "01101110011101100110111110001111",
        1614 => "10011000011100100111000001110010",
        1613 => "01110000011100110111001001100100",
        1612 => "10000001100110110111010010001011",
        1611 => "10001001100011101000100110010001",
        1610 => "01110101011101111000100001100010",
        1609 => "01100111011001100110011001101101",
        1608 => "01110010100000010111000010001010",
        1607 => "10010100011101010111000001110111",
        1606 => "01110010011100100111000101011000",
        1605 => "01101100101011111000000010101001",
        1604 => "10001111011111111000100010010110",
        1603 => "10100010100110010110100101101010",
        1602 => "01100100011100111000001010001100",
        1601 => "10011000100100011000101110101001",
        1600 => "10000101011101010111011101110010",
        1599 => "01110001011100010110111101011110",
        1598 => "01100010101010001000001101111110",
        1597 => "10000100100111110111111010001000",
        1596 => "01111010100000101000000110000101",
        1595 => "01111001100011110110110101110001",
        1594 => "01111001011101010111111110010101",
        1593 => "01111011011100110111010001110110",
        1592 => "01110001011101010110111101110000",
        1591 => "01110011011011100110100001111111",
        1590 => "10001000011010101000101101111000",
        1589 => "10000111100101100111000110001010",
        1588 => "01110101011101111000011010010010",
        1587 => "10001010100010011001101010001010",
        1586 => "10000000011101010111101001110011",
        1585 => "01110010011101110111010101110011",
        1584 => "01111001011110111000110110000101",
        1583 => "01101000101001010111000110001100",
        1582 => "10000101011101101010000101110111",
        1581 => "10000111100101111001011110000010",
        1580 => "01111001100010011000001010000001",
        1579 => "10000100011101010111010001110001",
        1578 => "01110010011110000111010001101110",
        1577 => "01101111011101100111010101110110",
        1576 => "10011111011111000111001110100011",
        1575 => "10000110011111001000100010010000",
        1574 => "10010001100010101000011101111111",
        1573 => "10001110100101011001101010010000",
        1572 => "01111101011110010111100101110101",
        1571 => "01110001011101100111001001101111",
        1570 => "01100100011101000111010101110110",
        1569 => "10010001101010101000100010111111",
        1568 => "10011111100110101010100010101100",
        1567 => "10101001101001011000111110010100",
        1566 => "10001011100010111000110101111001",
        1565 => "01110111011100010111010101111000",
        1564 => "01110100011101000111011101110111",
        1563 => "01110000011010100111000110011101",
        1562 => "10010010100100111001100110011001",
        1561 => "10011000101100111000110010101000",
        1560 => "10011110100100001000000110001100",
        1559 => "10000001100000101000010001110111",
        1558 => "01110001011110010111001001110010",
        1557 => "01110111011100100111010101110010",
        1556 => "01110101011101010111000101111000",
        1555 => "01110001011011110111000001110000",
        1554 => "01101101011100100111010101111101",
        1553 => "01110111011100010111010101110100",
        1552 => "01110100011101100111100001110001",
        1551 => "01110001011100110111100001111000",
        1550 => "01110111011110000111100101110011",
        1549 => "01110111011101010111001001110001",
        1548 => "01110011011101110111000101110100",
        1547 => "01111001011100100111001101110010",
        1546 => "01110010011110010111001001110011",
        1545 => "01110110011110010111001001110011",
        1544 => "01110110011110100111100001111001",
        1543 => "01111000011100110111011001111001",
        1542 => "01110110011100110111100001110011",
        1541 => "01110111011101010111001001110100",
        1540 => "01111001011100110111100101110111",
        1539 => "01111001011101100111011001110001",
        1538 => "01110110011100100111001001110000",
        1537 => "01110101011101000111000101110100",
        1536 => "01010011000000000000000000000000",
        1476 => "01110101011100010111001001110111",
        1475 => "01110101011100000110110101110101",
        1474 => "01110101011011110111001001110011",
        1473 => "01101111011001100111011001101110",
        1472 => "01110010011100010111011001101111",
        1471 => "01110010011011110111100001111000",
        1470 => "01110100011101000111011101110100",
        1469 => "01111000011110000111000101110110",
        1468 => "01110101011010100110011001100110",
        1467 => "01011010010101000101100101011001",
        1466 => "01010111010011100101100101100011",
        1465 => "01011110010111100101110101100100",
        1464 => "01100111011100000111010101111010",
        1463 => "01110001011101000111010001110011",
        1462 => "01110011011101000111000001110001",
        1461 => "01110001011100000110010101101010",
        1460 => "01100010011100100111001001110011",
        1459 => "10000110100000101000001001110001",
        1458 => "01110111100001100111000101100101",
        1457 => "01100111011010110111001101111000",
        1456 => "01110111011101000111100101110111",
        1455 => "01110110011101010111100101110011",
        1454 => "01110011011110000111101101111000",
        1453 => "10000011011110010111010010001000",
        1452 => "01110010100000110111011101110000",
        1451 => "10110111011100111000101101111000",
        1450 => "01111011011110010111001101110000",
        1449 => "01110100011110000111011001110010",
        1448 => "01111000011110010111010101101111",
        1447 => "01100111011010101000100110001000",
        1446 => "10001011100100110111101010001100",
        1445 => "01110001011110110111000101101110",
        1444 => "01110001011101101000001110000011",
        1443 => "01111100011111000110101001110100",
        1442 => "01110001011110010111011101110010",
        1441 => "01110010011110000110111101101111",
        1440 => "01110001100000111001010001111001",
        1439 => "10011101011101110111111001101110",
        1438 => "01101011011011000111000001101000",
        1437 => "01101111011011110110110101110010",
        1436 => "01101101011010100110011101101101",
        1435 => "01110010011110100111100101111000",
        1434 => "01110111011110000110101101101101",
        1433 => "01110111011110110111111010000111",
        1432 => "10000010011101101000010001100111",
        1431 => "01111011011011010110011101110000",
        1430 => "01110110011100110111100110001101",
        1429 => "01101000011001000111010001101110",
        1428 => "01101111011101110111000101110001",
        1427 => "01111000011101100110100101100101",
        1426 => "01100001011010110111101001110011",
        1425 => "01110001011111101000101110001111",
        1424 => "01110111011100010110010001101111",
        1423 => "01110101011010100111000101101001",
        1422 => "01101010011100100110100001111001",
        1421 => "01111100011110000111010101110110",
        1420 => "01110010011100110110100001100101",
        1419 => "01011101010110011000000001101111",
        1418 => "01110001011101010110111001110110",
        1417 => "01110101100100000110101101011110",
        1416 => "01110111011010110110101001101100",
        1415 => "01111000100011101000100101110101",
        1414 => "01111110011100000111011001110010",
        1413 => "01110010011101010101110101100010",
        1412 => "01101110011000101000011110000011",
        1411 => "01110111011100010110101010010010",
        1410 => "10000000100001101001100010100010",
        1409 => "01110101011011001000110110001010",
        1408 => "10001000100001000111110101111010",
        1407 => "01101100011110000111001001110110",
        1406 => "01101111011011100101111101100001",
        1405 => "01110011011101001001000101111100",
        1404 => "01101011100110001000111110001111",
        1403 => "10001100101001000111111101110111",
        1402 => "01111110100001111000111010010010",
        1401 => "10001111011110100111010001101011",
        1400 => "01011100011101000111100101111001",
        1399 => "01110100011010000110100101100101",
        1398 => "01111010011110011000111110011100",
        1397 => "10000011100000111001001110001111",
        1396 => "10100011100011110111111010001010",
        1395 => "01111100011111111000011110010111",
        1394 => "10010111100000100111000101011010",
        1393 => "01101001011100010111011101110110",
        1392 => "01110000011100110110010101001000",
        1391 => "01111011100110100111010101110000",
        1390 => "10010001011111111010000110100001",
        1389 => "10001001100001000110011110001000",
        1388 => "10100001100011111001100010010000",
        1387 => "10010011100100101000010010001111",
        1386 => "01111110011110100111100101110100",
        1385 => "01111000011010000111001001101000",
        1384 => "01110011100011001000010010000110",
        1383 => "10100101100000001010001010010100",
        1382 => "10000111100000010110101110101111",
        1381 => "10010011100010011000011110000110",
        1380 => "10011000100100111010001010011111",
        1379 => "01101111011011000111011001111000",
        1378 => "01101111011101000111000101100100",
        1377 => "01110100100101001010010010011011",
        1376 => "01111111100011001000101010001101",
        1375 => "10100100011101100110110010101101",
        1374 => "10100100101000011001110010001100",
        1373 => "10011010100111101000100101110101",
        1372 => "01101000011011100111010101110110",
        1371 => "01110100011010110110110001110110",
        1370 => "01101111100011101010100110001100",
        1369 => "10001000011110110111100010001111",
        1368 => "10000110011001110111011011011101",
        1367 => "10011101101001110111110010101011",
        1366 => "10110000100100101000000101011111",
        1365 => "01100011011001100111001101111000",
        1364 => "01110101011100100110001101010101",
        1363 => "01011100011101000110111001110110",
        1362 => "01111101100000001000111110100011",
        1361 => "10100101010101100100110010110110",
        1360 => "01111011101101001010101110010001",
        1359 => "10001110100011111000000001100100",
        1358 => "01101111011011000110111101111001",
        1357 => "01110100011011110110011001101010",
        1356 => "01100011100001101000101101110111",
        1355 => "10010001011111110111111101100110",
        1354 => "01101111010100010110010110010001",
        1353 => "01111100011100111000100101111001",
        1352 => "01111001011011010110011101101000",
        1351 => "01101001011011110111001001111000",
        1350 => "01110001011100100111000001101101",
        1349 => "10000111011111101000100010000111",
        1348 => "01111011100011010111100110001001",
        1347 => "01101010010111010110111101101110",
        1346 => "01111011011011100111010101111111",
        1345 => "01111010011110000111111001101000",
        1344 => "01101100011101100111011001110010",
        1343 => "01110110011100001000111010001101",
        1342 => "10001011011010001000100101110110",
        1341 => "01110000100000000111001001100111",
        1340 => "01101010011001010110100001101011",
        1339 => "01111111011011111000100001110001",
        1338 => "10001010100001111001000001111001",
        1337 => "01110101011111000111010101110010",
        1336 => "01110110011110110111101110001100",
        1335 => "10011011100011101000010001111111",
        1334 => "01111101011100110111011101100101",
        1333 => "01100111011000100110100001100011",
        1332 => "01110100011011101000001101111110",
        1331 => "10000110100001001001000110000010",
        1330 => "01110011011100100111000001110010",
        1329 => "01111001011110100111000101111101",
        1328 => "10011101100000000111001101110100",
        1327 => "01110100011010000110111001100111",
        1326 => "01100000011001110110100001101111",
        1325 => "01110010011100101000100001111101",
        1324 => "01111100011111001000110001111101",
        1323 => "01101110011100100111100001111000",
        1322 => "01110100011011100111001101111101",
        1321 => "10011001100010100111110110000011",
        1320 => "10001011100010010111111110001011",
        1319 => "01111101011111010110100110010000",
        1318 => "10000111011110111000001001111000",
        1317 => "01110100011100000111110001111110",
        1316 => "01111001011110000111001001110011",
        1315 => "01111001011100100111011010001110",
        1314 => "10010010100111111001111110011101",
        1313 => "10010011011101111000000010000010",
        1312 => "01110100011101010111110101110100",
        1311 => "01101111011000110110011001100010",
        1310 => "01110001011001100111011101111000",
        1309 => "01111001011100100111010101110111",
        1308 => "01110001011101100111100101110001",
        1307 => "01110110011101010111001101110111",
        1306 => "01110010011001100110100101100001",
        1305 => "01100000010110010011111001001110",
        1304 => "01011000010110100101010001010111",
        1303 => "01101011011011110111011101110011",
        1302 => "01110100011100110111001101110011",
        1301 => "01110001011100010111100101111000",
        1300 => "01101111011011100110111001101100",
        1299 => "01101111011010100110111001100100",
        1298 => "01100101011010100110001101011000",
        1297 => "01011110010111100110101101100110",
        1296 => "01100110011100000111100001110110",
        1295 => "01110110011110010111010001110010",
        1294 => "01111001011100100111011101111001",
        1293 => "01110101011100000111000101110011",
        1292 => "01110101011100100110111101101000",
        1291 => "01100011011101010110110101100011",
        1290 => "01101001011100100111001101101100",
        1289 => "01100111011011100111010101110110",
        1288 => "01110001011101100111100101110100",
        1287 => "01110001011101010111011101111010",
        1286 => "01110100011101000111100001111001",
        1285 => "01111000011100010111010101110001",
        1284 => "01111000011101010111000101111000",
        1283 => "01110111011110010111001101110011",
        1282 => "01110110011110010111100101111000",
        1281 => "01111001011101000111001001110011",
        1280 => "10001001000000000000000000000000",
        1220 => "01110010011100010111010101110010",
        1219 => "01110011011101100111011101110100",
        1218 => "01110100011101010111011101110010",
        1217 => "01110010011100110111000101111001",
        1216 => "01110010011101100111000101110010",
        1215 => "01110110011101000111010001110001",
        1214 => "01110110011110010111001101110111",
        1213 => "01110101011101010111001001110111",
        1212 => "01110111011100110111011101111010",
        1211 => "01110010011010010111000001111011",
        1210 => "10001011011111010111111110001100",
        1209 => "10000001011101010110100001100101",
        1208 => "01100111011011010111011001110110",
        1207 => "01110111011110010111011101110101",
        1206 => "01110001011101000111011110000001",
        1205 => "10001011100011011000111010000001",
        1204 => "10001100100101011010000110101111",
        1203 => "10111000011111111011000110101010",
        1202 => "10101011100111101001111001111000",
        1201 => "01111001011111010111010110000001",
        1200 => "01111001011110010111011001110101",
        1199 => "01110100011110100111000101111010",
        1198 => "01111111100010110111011010001001",
        1197 => "10000001101000101010110110000000",
        1196 => "10100001101000011010011110001101",
        1195 => "10001011100001111010011110001010",
        1194 => "01111011011111000111110101111011",
        1193 => "01111001011101010111011001110100",
        1192 => "01110011011101000111100010000000",
        1191 => "10000101100000000111100110001101",
        1190 => "01110111011011110111011110001011",
        1189 => "01110010100000110111001010000110",
        1188 => "10000001101001000111011110011001",
        1187 => "01101101100001111001000010000111",
        1186 => "01111111011110000111011101111000",
        1185 => "01110110011101001000000010001011",
        1184 => "10010010100010110111101110000101",
        1183 => "10001101100110100111011110000111",
        1182 => "01111110100010001000000010000000",
        1181 => "01111110011100010111111101111011",
        1180 => "10000011011100010110110110010100",
        1179 => "01111010011100100111100001111001",
        1178 => "01110100011101000111110010000100",
        1177 => "10000111100110111001101010011110",
        1176 => "01111110100000001000110001110010",
        1175 => "01111110100000100111101001111100",
        1174 => "10001011011111101000010010001001",
        1173 => "10100100100100100111101110010000",
        1172 => "01111001011100000111001101110100",
        1171 => "01111001011100111000000001111100",
        1170 => "10000111101011000111110001111111",
        1169 => "10010110100010011000111110001011",
        1168 => "01110101011100111000100001111000",
        1167 => "10001010100000001010000110010110",
        1166 => "01111000100100011010011101111111",
        1165 => "10000010100000000111010101111000",
        1164 => "01110100011100010111000110001001",
        1163 => "10010101100000101001001010011100",
        1162 => "01110011100010000111001001110000",
        1161 => "01111101011011101000100110000000",
        1160 => "10000110100011100111010010101000",
        1159 => "01110110100110100111010010100101",
        1158 => "01111100011111100111010101110110",
        1157 => "01110110011011110110100110001110",
        1156 => "10010000100011000111011101110001",
        1155 => "10000001011010011000100101111111",
        1154 => "01111111011111110111100101110011",
        1153 => "01111110011110110111010101110101",
        1152 => "10010010101101101001000110100111",
        1151 => "01111011011101110111100001111001",
        1150 => "01110101011100000110010001111010",
        1149 => "10001100011100001000010001111111",
        1148 => "01111111100110101001000101111111",
        1147 => "01111000011010010110100001100111",
        1146 => "01110001011101010111011101110100",
        1145 => "01101101101001111000100101111101",
        1144 => "01111010011010110111001001111001",
        1143 => "01110000011010110110101101111101",
        1142 => "10001111101001010111100110011001",
        1141 => "10000000011001100111100101101000",
        1140 => "01111010011011110111101101111011",
        1139 => "01110110100000000110100001110000",
        1138 => "01101000011011110111001001101111",
        1137 => "01110100011100110111011101110101",
        1136 => "01101110011011010110011010010010",
        1135 => "10001101011001011000100101110111",
        1134 => "01111001100111010111000101111010",
        1133 => "01101101011011100111110010001110",
        1132 => "10000010100001111000111001111001",
        1131 => "01101111011110110110111101110011",
        1130 => "01101111011100110111100101111000",
        1129 => "01110100011100100101100101110111",
        1128 => "01110100100010100111000101111100",
        1127 => "01100111011010010110100101110000",
        1126 => "01110111011111010111111010001010",
        1125 => "10000001100110011000000010000000",
        1124 => "10000001011101010111001110000000",
        1123 => "01110101011101010111001001110111",
        1122 => "01110011011100110101111100111000",
        1121 => "01011001011011010110111110000111",
        1120 => "10000011011100110111001001100101",
        1119 => "01101011011101111001101010101000",
        1118 => "10010110100000010111111101111010",
        1117 => "10100001011100101001011110000100",
        1116 => "01110010011101000111010101110001",
        1115 => "01110101100011000111010100101011",
        1114 => "00111110010101000101111101101111",
        1113 => "01100111011010010110010001101100",
        1112 => "10001000011101001001011110001111",
        1111 => "10001110101000010111110110000100",
        1110 => "10001110101001010111010101110111",
        1109 => "01101100011101110111011101110100",
        1108 => "01110001100010111101001011000101",
        1107 => "01110011010111000110100001100111",
        1106 => "01101001011100100110111101110100",
        1105 => "01110010100001101010111010001011",
        1104 => "10001011100001001000100110010010",
        1103 => "10010000100101100111011001110100",
        1102 => "01100010011101000111100101111010",
        1101 => "01111010100101011110000011110011",
        1100 => "10111110011010010111001001110000",
        1099 => "01101111011010100110100001101101",
        1098 => "01110100011110101000011010011000",
        1097 => "10000110100101011010000110011100",
        1096 => "10010100011011100111001001110000",
        1095 => "01100111011101000111011101111000",
        1094 => "01110111100010111011101111010111",
        1093 => "10011000100111111011011001110101",
        1092 => "01110101100000110111100101100111",
        1091 => "01100110011100000111001001111111",
        1090 => "10010001011111100110110001111100",
        1089 => "01110100100000010110111001010100",
        1088 => "01100010011100000111001001110011",
        1087 => "01110101100010001011001111000110",
        1086 => "10110001011100111000100010010111",
        1085 => "10001100011110011000000001111110",
        1084 => "01110000011100110111001101111000",
        1083 => "10000000100000111000100101111110",
        1082 => "01101101011110100110101001000010",
        1081 => "01100101011110000111000101110111",
        1080 => "01111000011111101010110010101011",
        1079 => "10010111100101011000100001111110",
        1078 => "01110101100000110111110110000011",
        1077 => "01100100100001110110101010000010",
        1076 => "01111101100101100111010010110001",
        1075 => "01111001011111000110110001001110",
        1074 => "01101000011101010111100101110110",
        1073 => "01110110100001001001011110100101",
        1072 => "10001011100011110111000110001001",
        1071 => "10011010100000010111110101110111",
        1070 => "01111000100010110111100010000101",
        1069 => "01111000011101100111011001111001",
        1068 => "01110111011101010111001001100000",
        1067 => "01100110011110010111100101111000",
        1066 => "01110010011111011001001010010100",
        1065 => "10001100100011100111101010100100",
        1064 => "01110100100001011001000110000011",
        1063 => "01101100011101011000001001111111",
        1062 => "10001000100111110111011001110011",
        1061 => "01110100011000100110001001011111",
        1060 => "01101111011101000111011001111001",
        1059 => "01110011011110001000101110011100",
        1058 => "10001110100000011001011101101011",
        1057 => "10001011101111101001001010000000",
        1056 => "11010111011110000111000110100111",
        1055 => "10101001011101010110111101100111",
        1054 => "01101110011001010110000101101101",
        1053 => "01110010011100100111100001110111",
        1052 => "01111001011110100111110001111110",
        1051 => "01110001100001011001100010010011",
        1050 => "10001000100110001000101001110100",
        1049 => "10001111011110100111110101111011",
        1048 => "01101101011100000111010001101111",
        1047 => "01110010011101100110101101110101",
        1046 => "01110110011101110111011101110001",
        1045 => "01110011011101010111011001101111",
        1044 => "01110010011100010110110001101110",
        1043 => "01110111011111100111111001110101",
        1042 => "01110000011010110110101001101101",
        1041 => "01101011011011000111001101110111",
        1040 => "01110110011100110111010101111010",
        1039 => "01110100011100110111000101111001",
        1038 => "01111010011101100111001001110001",
        1037 => "01111000011110000111100001110011",
        1036 => "01110001011100100111100001111001",
        1035 => "01110110011101100111010001110010",
        1034 => "01110010011100010111100001110001",
        1033 => "01110001011101100111001001111001",
        1032 => "01110100011101110111011101110111",
        1031 => "01110111011100100111011101111000",
        1030 => "01110011011101000111001001110100",
        1029 => "01110101011101110111010001110010",
        1028 => "01110100011101000111011101110010",
        1027 => "01110010011101000111001101110010",
        1026 => "01110101011100010111100101110111",
        1025 => "01110101011100010111000001110010",
        1024 => "11111110000000000000000000000000",
        964 => "01110111011110010111000101110011",
        963 => "01110010011100100111010001110100",
        962 => "01110011011101100111001101110011",
        961 => "01111000011101000111010001111000",
        960 => "01110111011101110111000101110101",
        959 => "01110100011101110111100001111001",
        958 => "01110110011100100111000101110010",
        957 => "01110010011110000111000001110001",
        956 => "01110001011101000111001001111001",
        955 => "01110001011101100111100001111001",
        954 => "01110011011101110111001101110010",
        953 => "01111000011100010111010001110010",
        952 => "01110010011101100111001101110010",
        951 => "01111001011110010111010101110011",
        950 => "01111000011100010111011001110000",
        949 => "01110011011101010111100101110011",
        948 => "01101111011100110111001101101111",
        947 => "01101010011100000110110101110111",
        946 => "01110101011100100111001101110101",
        945 => "01110010011101110111000101110110",
        944 => "01110110011100100111010101110010",
        943 => "01110101011100100111100001110010",
        942 => "01110010011100100111000101110000",
        941 => "01101101011101010111100101111011",
        940 => "01101111011010000110001101100101",
        939 => "01011000011000000110010001101010",
        938 => "01110010011101000111001101111001",
        937 => "01110001011101000111100001110111",
        936 => "01110001011110010111001001101101",
        935 => "01101101011011100111011010000001",
        934 => "10010010100101010111011101110100",
        933 => "01110101011110110111010001110110",
        932 => "01101111011010010111000001101010",
        931 => "01100111011010110111001101110001",
        930 => "01111000011101110111011101110000",
        929 => "01111001011101100111100001100110",
        928 => "01100100011010011000011110001100",
        927 => "01111111011110110111011010000101",
        926 => "10100111011010011001001010010001",
        925 => "01101010100111101000011001111111",
        924 => "01110101010111100110011101101011",
        923 => "01110101011100110111100001110110",
        922 => "01110111011101010110111001110000",
        921 => "01101110100000110111001010010111",
        920 => "10001111101000111001111110001000",
        919 => "10001001100110111001010110100101",
        918 => "10001100100011001000101110100111",
        917 => "01111100011010100110011001101000",
        916 => "01110101011100100111010101110101",
        915 => "01110110011101000110110101101101",
        914 => "10000000011110001001000110011010",
        913 => "01111100100101001000001110001000",
        912 => "10001110101000110111111110011111",
        911 => "10010100101001101001111101101110",
        910 => "10011101011101010111010001101110",
        909 => "01110011011101010111100001110111",
        908 => "01110011011100100110100001110011",
        907 => "10001101100111001000100001111111",
        906 => "10000101100001001000101110000011",
        905 => "10001011100110011000011110100011",
        904 => "10101010101000011001110001111000",
        903 => "10001001100100010111100101110011",
        902 => "01110010011110100111010101110110",
        901 => "01110101011100101000001110000100",
        900 => "10001001011101110111110101111010",
        899 => "01111001100011001000101110001111",
        898 => "01111001011101001001101010110000",
        897 => "01111101100011111001000110001001",
        896 => "10011110100000000111001001100000",
        895 => "01110011011101100111001001110010",
        894 => "01110101011010111000101010000110",
        893 => "10000111100010111000010110000011",
        892 => "10000110100000001000100001110101",
        891 => "01110111100100001000100110000101",
        890 => "10101100101011011001111110010110",
        889 => "10001000100001011000001101011000",
        888 => "01110000011101110111100001111000",
        887 => "01101111011000111000100010000001",
        886 => "01111000100001001000100101111011",
        885 => "10001010100010100111001010000001",
        884 => "01111101100010000111100001111001",
        883 => "10110100100100011001110010001110",
        882 => "10010110101001011000010101011011",
        881 => "01101000011101010111011101110100",
        880 => "01110111011000111000110010000110",
        879 => "10000001011110111000110110000110",
        878 => "01111010011110101000001001111011",
        877 => "01111011100101111000101110010101",
        876 => "10010001100010010111111110010001",
        875 => "10010000100100000111000001011001",
        874 => "01110001011110100111001001111000",
        873 => "01110001011001100111111010010000",
        872 => "10010001100011111000101001111001",
        871 => "01111101011110000110010110001101",
        870 => "01111111011100110111100110001011",
        869 => "10100100100101101000111110001101",
        868 => "01111010100100101000101001011110",
        867 => "01110010011100010111011101110101",
        866 => "01110010010110100101100110011001",
        865 => "10110101100011101001011101111010",
        864 => "10000100011100100110110001111101",
        863 => "10000100011011111001011010010000",
        862 => "01111001100011110111100101110110",
        861 => "10001001101010011000100101110001",
        860 => "01101111011101010111000101110010",
        859 => "01110001010110000110000110011001",
        858 => "10111101101001011001001001111001",
        857 => "01100011011011010111010001111100",
        856 => "01101010011011111001001010010001",
        855 => "10100001100001111000111010010011",
        854 => "10100010100011010111110001110011",
        853 => "01101011011101100111011101110000",
        852 => "01110100010110000101001001111000",
        851 => "10011011011011101000010101111001",
        850 => "01111010011001110110011101110101",
        849 => "01011100011101001001011110010001",
        848 => "01110111100000101001101110000110",
        847 => "10010110011101000111110001110101",
        846 => "01110010011100100111100101110100",
        845 => "01110011011001100101100001110001",
        844 => "01110100011001000111000101110010",
        843 => "01101000011001010110011101100100",
        842 => "01011100011001110111010001101101",
        841 => "01101110011101110110111110000000",
        840 => "01111111011100010110110001110010",
        839 => "01101011011100110111001101110100",
        838 => "01110000011001010101101101101000",
        837 => "01101101011011010111101001101110",
        836 => "01100100010110100101100101011101",
        835 => "01100111011011110101110001101100",
        834 => "01110000011001010110101101110000",
        833 => "01111100011011100110100110000010",
        832 => "01110100011100110111101001111001",
        831 => "01101111011011000110010101100001",
        830 => "01100101011011010111000101101010",
        829 => "01100000010110100110110001101000",
        828 => "01011100011000000111010001101001",
        827 => "01101111011100000111100001110010",
        826 => "01110000011011100111010001110111",
        825 => "01101101011101010111010101110101",
        824 => "01110101011100110111000010001000",
        823 => "01110101011011100111010001101001",
        822 => "01101000011010000110101101100111",
        821 => "01110001011100110110001101110001",
        820 => "01111010011100000111010101110011",
        819 => "01111111011000100111011001110011",
        818 => "01101111011110000111000101111001",
        817 => "01110110011110110111010110001110",
        816 => "10001000011100100111010101101111",
        815 => "01101000011001100110111101101010",
        814 => "01110110011010000110011101110000",
        813 => "01101110011010000111010101110111",
        812 => "01110101011000110110110001110101",
        811 => "01101111011110000111010001111000",
        810 => "01111010011101110111001001111111",
        809 => "10011110011100101000101010000110",
        808 => "10011010100011011000010001110011",
        807 => "01101101100000010110110001110101",
        806 => "01101011100011110111101110000110",
        805 => "01101100011100100110100001110110",
        804 => "01101111011100100111010101110110",
        803 => "01111010011110000110101101100000",
        802 => "10001011100011001000011110000101",
        801 => "10000000100000011001000110010011",
        800 => "10000010100001011000001101111111",
        799 => "01111101100001110111000110000001",
        798 => "01110101011111010111100001111011",
        797 => "01110100011110010111001001110111",
        796 => "01110011011101010110110010000001",
        795 => "10001101100001100111111101111001",
        794 => "10001101100010000111110110000011",
        793 => "10001100100011001001000010001100",
        792 => "10010000100011111001000110001000",
        791 => "10000111100000010111010001110110",
        790 => "01111000011100110111010001110010",
        789 => "01110111011110000111000101110110",
        788 => "01111110100001101000111110000111",
        787 => "10001100100001001000010110000011",
        786 => "10000011100010111000101010010011",
        785 => "10010100100100111000100110001111",
        784 => "10001100011111100111001001111010",
        783 => "01110111011100000111000001111001",
        782 => "01110111011100100111001001111001",
        781 => "01111100011110100111101001111000",
        780 => "01111110011111000111011101110101",
        779 => "01111000011110001000001010000111",
        778 => "01111011011110100111110010000000",
        777 => "01111111011111010111100001111001",
        776 => "01110001011110010111001101111000",
        775 => "01110111011101010111001001110100",
        774 => "01111001011110010111000101110110",
        773 => "01110100011110010111010101110110",
        772 => "01110011011100110111001001111001",
        771 => "01110101011100010111000001110110",
        770 => "01110010011100100111011001110101",
        769 => "01110011011101000111001001110101",
        768 => "01101111000000000000000000000000",
        708 => "01111001011100110111001101110110",
        707 => "01110100100000001000000001111011",
        706 => "10000011100001001000000101111111",
        705 => "01111100100000011000011001111011",
        704 => "01111001011111000111010101111000",
        703 => "01110011011101110111000101110010",
        702 => "01110111011110100111011001110011",
        701 => "01110001011110010111011001110000",
        700 => "01110100100000100111100001110110",
        699 => "10010110100101101001011110001100",
        698 => "10011101100101011001010110000001",
        697 => "10000101100011011000110010000100",
        696 => "01111011011000100110100001101111",
        695 => "01111001011110000111100101110110",
        694 => "01110001011110000111011101110001",
        693 => "01110001011101010111010101110000",
        692 => "01111111100100011001000010011000",
        691 => "10011010101000001001100010101110",
        690 => "10110110100101111010000110010100",
        689 => "10000100011100110111011010000100",
        688 => "01110111011101010111010001110111",
        687 => "01110100011101100110111101101110",
        686 => "01011011011001010110100001101011",
        685 => "01101101011010001000010101110011",
        684 => "01111001011110111000111101110000",
        683 => "01111101100000010111010110001011",
        682 => "10001110100101111001101101111111",
        681 => "01110111011101010111001101110101",
        680 => "01110001011100010111010001101111",
        679 => "01010110010101000101000101011001",
        678 => "01101000011011010111001001110000",
        677 => "01111010011011100110001001100100",
        676 => "01100111011011100110111001011101",
        675 => "10011100100011110111101001110010",
        674 => "01100011011100110111011001111001",
        673 => "01110001011100110111010101101111",
        672 => "01011001010100010101011101100011",
        671 => "01110101011010110110101001110111",
        670 => "01110000011101110110000001111101",
        669 => "01100111011101010111001001110111",
        668 => "10000001011100010111000101011110",
        667 => "01100010011010010111010101111010",
        666 => "01110110011100110111000001110100",
        665 => "01010111010100000101101001100101",
        664 => "01100110011010000110100101110100",
        663 => "01101000010111110110010001110001",
        662 => "01101111011101010110111101110100",
        661 => "01011101010111010110001101011010",
        660 => "01101000011100000111010101110100",
        659 => "01110100011101010110110001101110",
        658 => "01100010010100010101111001011010",
        657 => "01100111010110100110000101100000",
        656 => "01100110011110110111010001111011",
        655 => "01101110011011100110111001110011",
        654 => "01100110010110110110001001011110",
        653 => "01100110011100010111010001110001",
        652 => "01110111011110010111010101101111",
        651 => "01010101010110100110111001110001",
        650 => "01110010011001000110101001101000",
        649 => "01101000011111100110111001110100",
        648 => "01110001011000000111001101110011",
        647 => "01100111011011000110111101110100",
        646 => "01101101011111000111011001110110",
        645 => "01111001011101010111011101101101",
        644 => "01011101011101011000000001110011",
        643 => "01110100011101100111011101110010",
        642 => "01110001011100101000001101101110",
        641 => "01111000011101000110111101101110",
        640 => "01101100011001110111111101111101",
        639 => "01101110011101110111010001110001",
        638 => "01110000011101110111110110000010",
        637 => "01110110100000000111010110001100",
        636 => "01101110100011010111011001110111",
        635 => "10001000100001011000000110000110",
        634 => "01101101011001110111001001110100",
        633 => "01101111011101011000000010000010",
        632 => "01101010011100010111011001110001",
        631 => "01110001011011110110011101101000",
        630 => "01110010011100101001010110011000",
        629 => "10010010011110111001100001111000",
        628 => "10001011010110010111110101101110",
        627 => "01011010011010000111000001111001",
        626 => "10100111011101110110111001111101",
        625 => "01101101011101110111001101110100",
        624 => "01110010011011100110000001101011",
        623 => "10010111101000011000111110010110",
        622 => "01111011101000111100000001011111",
        621 => "10001100011001100110110001011100",
        620 => "01100111011100010110101101101100",
        619 => "01110001011110100111001101110000",
        618 => "10000011011101110111000001110110",
        617 => "01110010011110000110111001110010",
        616 => "10010100100010100111000110011111",
        615 => "11000011100011011000100110001001",
        614 => "01110001011100010110001001011001",
        613 => "01100011011101000111000101111010",
        612 => "01110110011101101001000110001001",
        611 => "10001001100000000111101001110100",
        610 => "01110011011101010111110001111010",
        609 => "01101100011110011010000010010000",
        608 => "01100111011100110111101010001110",
        607 => "01111010011100010101100101001111",
        606 => "01110000100001100111000001101000",
        605 => "10000000101100101000001110001110",
        604 => "10011000100010100111011001111000",
        603 => "01110011011111010111011001100101",
        602 => "01101110101010111000111001111001",
        601 => "01111010101000001001011110100111",
        600 => "10101011011011010101000001011101",
        599 => "10011000011100010111000011011010",
        598 => "10101001011110011000100010011110",
        597 => "10100000100110010111111001110101",
        596 => "01110111011100110110111001100101",
        595 => "01110000100111001001001010101010",
        594 => "10000010101010011000111110001011",
        593 => "10100110101100111000100010000110",
        592 => "10010100101101101001000001101110",
        591 => "10010001100001100111111010001101",
        590 => "10010001100110110111110001110101",
        589 => "01110010011110110111011101101011",
        588 => "01110111100111001001101010101011",
        587 => "10100001100010111000011010110100",
        586 => "10001100100010001001100001100111",
        585 => "01100110011101101001000101111000",
        584 => "10000110100011101000110110001111",
        583 => "10010001100010110111111101110010",
        582 => "10000000011101010111100001111100",
        581 => "10000011100100011001011101110110",
        580 => "10010100100101111011010110001111",
        579 => "10010100101010010111100110100011",
        578 => "10000010011110001000110010000111",
        577 => "10000110100100111000101010010001",
        576 => "10001111100000000111110101110111",
        575 => "01110101011101100110101001110010",
        574 => "10001100100100100111010110010101",
        573 => "10000010100111101000001010001000",
        572 => "10011000100010100110111110011100",
        571 => "10010010011111111001000110011000",
        570 => "10100101100011101000101110001100",
        569 => "10010101100000000111101001110010",
        568 => "01110100011110010111001001111000",
        567 => "10000000100000111000110110100100",
        566 => "01110111101000111000101010001011",
        565 => "10001001011011011000110110001111",
        564 => "01111011100011101000110101111011",
        563 => "10011001100011000111110110001010",
        562 => "10010011011111110111010101111001",
        561 => "01111000011110000111000101101101",
        560 => "01100101011101001000011101110011",
        559 => "01111001011111111000101010000101",
        558 => "01111100011110110111010010010010",
        557 => "10101110100011101000111010011010",
        556 => "10010000100101011000110101111111",
        555 => "10000110011101000111010001110101",
        554 => "01110111011110000111000101110000",
        553 => "01101111011010010110011101011011",
        552 => "01100101011011100110111001110011",
        551 => "01110001011100101000000110001011",
        550 => "01110111011101101001010110010010",
        549 => "10000100011110100111110001110010",
        548 => "01110100011101000111100101110010",
        547 => "01110101011101100111011101110001",
        546 => "01110100011100010111010101101111",
        545 => "01101010011010110110011101100110",
        544 => "01100101011001010110100001100100",
        543 => "01011100010101110101111101101001",
        542 => "01101011011011000111010001110110",
        541 => "01110001011100100111001101110101",
        540 => "01110111011100110111100101110111",
        539 => "01110111011110000111011001110111",
        538 => "01110100011101110110111001110001",
        537 => "01101101011011110110100101101011",
        536 => "01101001011010000111001101110010",
        535 => "01110101011101110111101001111000",
        534 => "01110100011100010111001101111001",
        533 => "01110011011101100111001101110101",
        532 => "01110000011110010111001001110001",
        531 => "01110010011101100111001001110101",
        530 => "01110100011100010111010001110101",
        529 => "01110100011100000111000001110111",
        528 => "01110101011101110111010001111000",
        527 => "01110101011101010111000101111000",
        526 => "01110001011110010111100001110001",
        525 => "01110001011100110111000101110111",
        524 => "01110100011110010111011001110110",
        523 => "01110100011110000111000101110100",
        522 => "01110111011101110111101001111001",
        521 => "01110001011101100111000101111001",
        520 => "01111001011101110111100101110011",
        519 => "01110011011110010111001001110110",
        518 => "01110110011101000111000101110010",
        517 => "01110000011101110111001001110001",
        516 => "01110111011110000111011101110101",
        515 => "01110100011100110111001001110001",
        514 => "01110101011110010111000101110100",
        513 => "01111001011101000111001101111001",
        512 => "11010100000000000000000000000000",
        452 => "01111001011110010111100001110111",
        451 => "01110011011101100111000101110011",
        450 => "01110101011110010111001101110101",
        449 => "01110001011101100111100101110101",
        448 => "01111001011101010111100001110100",
        447 => "01111010011101110111010001110011",
        446 => "01110010011110000111101001110011",
        445 => "01110110011101100111010001110110",
        444 => "01110001011101000111000001101010",
        443 => "01101111011100010111000101101010",
        442 => "01100111011010110111010001110100",
        441 => "01110011011011000111000101110100",
        440 => "01110101011010110111010101110111",
        439 => "01110110011101110111100001110011",
        438 => "01110100011101100111100101110100",
        437 => "01101101011100110110111101111011",
        436 => "10001001100001011010101110100000",
        435 => "10100110101001100111110010001101",
        434 => "10101011101001000111000101110000",
        433 => "01110001011100000110001001101101",
        432 => "01111001011100110111100101110011",
        431 => "01110001011100100111010101101100",
        430 => "01110001011100000111001010001000",
        429 => "10111111100111100110011111001000",
        428 => "10001010101010001001001010010101",
        427 => "10100011011111011000001110011111",
        426 => "01110000011001100101110001100110",
        425 => "01101011011101100111011101110110",
        424 => "01110101011101010111001001101110",
        423 => "10000100100000001000000110001000",
        422 => "10010101101000010111101010000110",
        421 => "10000101011110111001011110000101",
        420 => "10000010011111000111111010011111",
        419 => "01101011011010000110101101110100",
        418 => "01110100011110010111011001111001",
        417 => "01110111011100100111000001101110",
        416 => "01111101011110111000101001101011",
        415 => "01110100011111110111110001110100",
        414 => "01111111100001010111100101111101",
        413 => "10000011011110100111100001101110",
        412 => "10001010100011010111100001111101",
        411 => "01110101011100010111001101110001",
        410 => "01110100011101100110111101100010",
        409 => "01110110100011110110111110001110",
        408 => "01111111011111101001000101110010",
        407 => "01110011011101111000001001101000",
        406 => "01111101011010111001010101110110",
        405 => "10100011101000000111010001110110",
        404 => "01101010011101100111011001110101",
        403 => "01110111011101100110100101100111",
        402 => "10001010100011001011000110011101",
        401 => "10001010011110000111100101101010",
        400 => "10000010011001011000001001111110",
        399 => "01110101100100100111110010001000",
        398 => "10101001011110010111011001101111",
        397 => "01100110011100010111001101111000",
        396 => "01110110011100100110010001101011",
        395 => "10100110101000100110101101110100",
        394 => "10000000100010001000001101111110",
        393 => "01110010011100100111001110000011",
        392 => "01110011100011101000111010000011",
        391 => "01101111100001101010010001101110",
        390 => "01100111011101000111001101110010",
        389 => "01111001011101000110001001110001",
        388 => "10010000011100110110111110000011",
        387 => "01110001011101100110110101110011",
        386 => "01110110011101011000010110001101",
        385 => "10010111100101101001001101111111",
        384 => "01110100100110000111010001101100",
        383 => "01101100011101000111010101110011",
        382 => "01111000011100000110001010000111",
        381 => "10001110011101010111101101110101",
        380 => "01110111011001100111011110000110",
        379 => "01110000100000111000100110010001",
        378 => "10001100100000111001110110001011",
        377 => "10110011011100000111000101110010",
        376 => "01110101011101100111010101110011",
        375 => "01110100011011110110100001101010",
        374 => "10000100011011000111000101101101",
        373 => "01100111011100111000100010001000",
        372 => "01111110100001101000101010011001",
        371 => "10000101100100100111110101110101",
        370 => "01110100011101010110101101101000",
        369 => "01111010011101010111001001110110",
        368 => "01110110011100000111101001100101",
        367 => "01101010011101000111001101110000",
        366 => "01111001100001000111011101111001",
        365 => "10000001100110101001000010001101",
        364 => "01111001011101011000011001110001",
        363 => "01110101011100110110011101101001",
        362 => "01110011011101100111010101111001",
        361 => "01110011011101010111101101100111",
        360 => "01100011011001110111010001101011",
        359 => "01111101011101001000001110000010",
        358 => "10000011100010101001100110001110",
        357 => "10011100100000010110100101101011",
        356 => "01101101011110010111100001100101",
        355 => "01110111011101000111011101110000",
        354 => "01111000011101010111110110010000",
        353 => "10011100100010000110101010101100",
        352 => "01110110011111010110111110001000",
        351 => "10011001011101111010100010011001",
        350 => "10010000011011101000000001111110",
        349 => "01111011100110001000001001110010",
        348 => "01111011011101110111100101110000",
        347 => "01110000011101110111100110111100",
        346 => "10110001101000011011000110001001",
        345 => "10011100011100111000011101111101",
        344 => "10000111100001101001111010001101",
        343 => "10000111011111001000110001101101",
        342 => "10100100011100001010010001111000",
        341 => "01111110011110010111011101110100",
        340 => "01110101100001100111100110010111",
        339 => "10010110100100010111100110000000",
        338 => "01110101011010010111000001111001",
        337 => "01111110101101001001101010001111",
        336 => "10001011100100101010001010100110",
        335 => "11000110100010101000111010000001",
        334 => "01110001011100010111011001110101",
        333 => "01110101011110100111001001110110",
        332 => "10010011100100001001001110010000",
        331 => "10011101100100110111011001101100",
        330 => "01011110011101010111100110011011",
        329 => "10000011100110001000100101111010",
        328 => "01110101100001000111010010010010",
        327 => "01101110011100110111011001110100",
        326 => "01110010100100001001011110011100",
        325 => "10011010100010011000111010000001",
        324 => "10000001011101101000101101111100",
        323 => "01100101011101110111110001101001",
        322 => "10000111011110001000101110010000",
        321 => "01111110100100110111011101110110",
        320 => "01110010011101100111010001110110",
        319 => "01111111100010011001000110110011",
        318 => "10001010100001011000111110000010",
        317 => "10010010100010110111011110001111",
        316 => "01110011011011101000101110000110",
        315 => "01111001100010101000101101110001",
        314 => "10011011100101101000100101111001",
        313 => "01111100011100110111010001110001",
        312 => "01110011011101100111111010011001",
        311 => "10101000011111001001010001110010",
        310 => "01110111100010000110111001111011",
        309 => "10001110011000000111110101101110",
        308 => "01101101100001000111001110100111",
        307 => "01101100011011100111010101110010",
        306 => "01110000011100010111011101110001",
        305 => "01110010011101111001001101110001",
        304 => "10011101011101010111011110000001",
        303 => "10011111011011111000110101111110",
        302 => "10001111100000001000000010011011",
        301 => "01110101011110101000001001111010",
        300 => "01110011011011110110111001101111",
        299 => "01110110011100100111011001110100",
        298 => "01111000011101101000111010000011",
        297 => "01101101011101110111111010010111",
        296 => "10001000011011011010000010000111",
        295 => "01111111100010011000000010010000",
        294 => "10100011011011011000011001110001",
        293 => "10000010011011000110101101110101",
        292 => "01110000011101100111100001110110",
        291 => "01111000011111001000010110000110",
        290 => "01111110100100001000000110100111",
        289 => "01110010101110011000101110110011",
        288 => "10100001110001010110010011011101",
        287 => "10001011100111001001000010000101",
        286 => "01110010011011000111000101110011",
        285 => "01110110011100100111010101110100",
        284 => "01111000011100010111010001110101",
        283 => "10000010100010000111110101110010",
        282 => "01110001100011101000001101110110",
        281 => "01110110011101010111100101110011",
        280 => "01110100011110010111010101111000",
        279 => "01110001011100100111001001110001",
        278 => "01110010011101010111100101110110",
        277 => "01110011011101000111001001111001",
        276 => "01110101011100110111001001110101",
        275 => "01110011011101010110111001101110",
        274 => "01110000011100110111000101110000",
        273 => "01110000011100000111100001110100",
        272 => "01110011011110010111000101110110",
        271 => "01110110011100100111010101110010",
        270 => "01110011011101110111010001111001",
        269 => "01110100011100010111011101110011",
        268 => "01111000011100010111010101110110",
        267 => "01110110011101110111100001110011",
        266 => "01110010011101000111100101111000",
        265 => "01111010011100100111100101110001",
        264 => "01111001011100100111011101111000",
        263 => "01110001011100100111001001110011",
        262 => "01110010011101000111011001111010",
        261 => "01110001011101010111100101111000",
        260 => "01110111011101000111011101110101",
        259 => "01110110011100000111001001110100",
        258 => "01110011011101000111001001111001",
        257 => "01111000011101100111000101110001",
        256 => "00000000000000000000000000000000",
        196 => "01110101011110000111100101110111",
        195 => "01111000011101100111100001111000",
        194 => "01110000011101000111001001110001",
        193 => "01111011011101100110100101111010",
        192 => "01110011011101110111011101111000",
        191 => "01111001011101100111001101111000",
        190 => "01110011011110100111100001110110",
        189 => "01111001011101010111010001110111",
        188 => "01111010011101111000100010001101",
        187 => "10001101101001001001011010011100",
        186 => "10010111101110001010010010101111",
        185 => "10100001101001011010110010100010",
        184 => "10100001100110101000111001111110",
        183 => "01110111011100110111001001110110",
        182 => "01110011011101000111011001101110",
        181 => "01111011011101101001001010011100",
        180 => "10001101100100101001010110011101",
        179 => "10010011101010101001100110100101",
        178 => "10100000101001011001001010011101",
        177 => "10010000100100001001110001110111",
        176 => "01110001011100010111011001111000",
        175 => "01110010011100100111000001101011",
        174 => "10001011100011111000011110001111",
        173 => "10001001100010001000101010000110",
        172 => "10000001011001110111000101110010",
        171 => "10000000100010110110101110010001",
        170 => "10000011011111000111100101110111",
        169 => "01110001011110010111011101110010",
        168 => "01110100011100010111010010000101",
        167 => "10000110100111001000101001111100",
        166 => "01111110011110000111001001110011",
        165 => "01101101011111110111000101101111",
        164 => "01110000011100100110100010000001",
        163 => "01101111011011000110100101100111",
        162 => "01110001011101000111000001110010",
        161 => "01110110011101100111011110000000",
        160 => "10000101011100100110110101111000",
        159 => "01101000011011110110111001101100",
        158 => "01011101011110010110100001111001",
        157 => "01110110100001110110111110001011",
        156 => "01110100011100100110011001101110",
        155 => "01110110011101100111101001111001",
        154 => "01110101011100110111010010000100",
        153 => "01110101011010000111011101110100",
        152 => "01110100011010110110100001110000",
        151 => "01100100010111000101111001100011",
        150 => "01100011011011010111000101110001",
        149 => "01110100011111100111100001101110",
        148 => "01101110011101110111000101110001",
        147 => "01111001011101110111101010000100",
        146 => "01110100011011110110100001110000",
        145 => "01111001011100010111100001110111",
        144 => "01100100011011000110101101011001",
        143 => "01011011011001110110110001110010",
        142 => "01101111011101010111111101101101",
        141 => "01100101011100100111000101110001",
        140 => "01110011011101000110110101101101",
        139 => "01100111011010010111000001111110",
        138 => "10000010011101000110011101110101",
        137 => "01100100011010000110110001110101",
        136 => "01101000011011100110111001111001",
        135 => "10001010011111010110100101100011",
        134 => "01101000011101000111001001110101",
        133 => "01110011011100010110110101010110",
        132 => "01011011011011010111010010000011",
        131 => "01101111011100100111111101111011",
        130 => "01111110100011010110101001101000",
        129 => "10010100101010010111000001110001",
        128 => "01111101100010010110011101100011",
        127 => "01101000011101000111011101110100",
        126 => "01110101011101100110110101011001",
        125 => "01100001011011110111010001110100",
        124 => "01110001011111101000000101111011",
        123 => "10010000011101111000010010000111",
        122 => "01110000100011000111100110010001",
        121 => "10001011011100000111000001100100",
        120 => "01101010011100100111100101110101",
        119 => "01111010011100110110010001010110",
        118 => "01100001100001000111000101111001",
        117 => "01101011100000111000111110001011",
        116 => "01111010011111000111001101110111",
        115 => "10001011100001110111000110001111",
        114 => "01111100011101001000001110000001",
        113 => "01110000011100000111001101110010",
        112 => "01110100011011100110110001010100",
        111 => "01100110011110110111000110000100",
        110 => "10001100100000001001110110001100",
        109 => "10001101011011100111101101110100",
        108 => "10001001100000110111101010001000",
        107 => "10000010100001000111111010000011",
        106 => "01110100011011000111100101111000",
        105 => "01110111011100010110100101010001",
        104 => "01011110011111101001010010010001",
        103 => "01111111100001101001010010001111",
        102 => "10001010011111001000111010000001",
        101 => "10000000100000110111110101110101",
        100 => "10000010101000010111111110010010",
        99 => "01110100011100000111011001110100",
        98 => "01110110011011000110000001010011",
        97 => "01101010100001111001110010011000",
        96 => "10011110100010001000101010011110",
        95 => "10010001100010011000111101111001",
        94 => "10000101100001000111100010001111",
        93 => "10100000011111111001001010110011",
        92 => "01101110011001110111001001111001",
        91 => "01110111011011110110101001100000",
        90 => "10100110101001101010101010001000",
        89 => "10010101100101011000110010001110",
        88 => "10010111100011001000010001110101",
        87 => "10010111100100111001011110010111",
        86 => "10011100101011011001100110001110",
        85 => "01100110011010000111000001111000",
        84 => "01110001011100110110100101100111",
        83 => "01110010101001011001110010111011",
        82 => "01111110100100001001110010010001",
        81 => "10011101100001001001010110011100",
        80 => "10010110101000011001011010110010",
        79 => "10010111100001010111111101101110",
        78 => "01100011011000000110110101110101",
        77 => "01111000011101010111001001100111",
        76 => "01110100011111010111100110000010",
        75 => "10001110100001010111011001111110",
        74 => "01101101011101110110011010000010",
        73 => "01111101100000101000010110001000",
        72 => "01110111101000000111011001101110",
        71 => "01101000011011010110111101111000",
        70 => "01110111011100110110111001110100",
        69 => "01110100100001100110110010001000",
        68 => "10000010100011011000101001111110",
        67 => "10011011100010100111110001111111",
        66 => "10000001100011100111111001111100",
        65 => "01110101101001000111011101100110",
        64 => "01100111011010100111001101110011",
        63 => "01110011011100010110111101111001",
        62 => "01111011011101111010110001101101",
        61 => "01111111100011000111111010001110",
        60 => "10000011100100001000010101100101",
        59 => "01110111011110010111100010101000",
        58 => "01100111011110010110111101100001",
        57 => "01100100011100000111011101110111",
        56 => "01110100011011010111000101101111",
        55 => "01111100011101010111010110001111",
        54 => "10000001100001101000101110011011",
        53 => "10011011100011111001100110010011",
        52 => "01111010011110100111100001110100",
        51 => "01101111011100000101101001100100",
        50 => "01101101011100100111000001110111",
        49 => "01110101011100000111000001101101",
        48 => "01101110011100010111011010010111",
        47 => "01110111101000101001000110010111",
        46 => "10001001100011111001101101111110",
        45 => "10011010011100001001010101110100",
        44 => "01101111011001110101111001101100",
        43 => "01110101011100110111001001111001",
        42 => "01110110011101010111001001101101",
        41 => "01101001011001110111000001110100",
        40 => "01110101011100100111001001101010",
        39 => "10001001011001111000111010001111",
        38 => "10111100011010010110111001101101",
        37 => "01101011011100000111010001111001",
        36 => "01110100011100110111010001110110",
        35 => "01110111011101010111001101110010",
        34 => "01110011011010110110011101101000",
        33 => "01100100011011100110111101101111",
        32 => "01110110011101000111000101101111",
        31 => "01101110011011000110110001101110",
        30 => "01110011011110000111010001110100",
        29 => "01110100011100110111100101110100",
        28 => "01110111011110010111011101110110",
        27 => "01110001011101010111000101110010",
        26 => "01110001011101000110111101101000",
        25 => "01100110011010100110011101101010",
        24 => "01101101011100100111001101110001",
        23 => "01110010011110010111000101111001",
        22 => "01110100011101110111011101110111",
        21 => "01110111011101110111011001110100",
        20 => "01110001011101000111001001110100",
        19 => "01110101011101010111001001110010",
        18 => "01110011011101010111000101110101",
        17 => "01110100011100010111001001110101",
        16 => "01110011011100100111100001111001",
        15 => "01111001011110000111100001111000",
        14 => "01110101011110010111011001110111",
        13 => "01110101011101010111011101110010",
        12 => "01110100011101010111100001110000",
        11 => "01110101011110000111100001110010",
        10 => "01110001011100110111010101110011",
        9 => "01110010011101010111100001110110",
        8 => "01110100011100010111001001110010",
        7 => "01110101011101110111000101110100",
        6 => "01110100011100100111010101110111",
        5 => "01111001011110100111100001110011",
        4 => "01111001011100110111100101110001",
        3 => "01110010011100100111011101110110",
        2 => "01110101011101000111011101110100",
        1 => "01110010011110010111010101110110",
        0 => "01100011000000000000000000000000",        
        -- here ends the generated array allocation

        others => "00000000000000000000000000000000"
    );

    signal rom_index: std_logic_vector (11 downto 0);
begin
    rom_index <= (in_rom_neuron_index & in_rom_input_index); -- combine the neuron and input index to adress the array
    out_weights <= rom_arr(to_integer(unsigned(rom_index)));
end RTL;
