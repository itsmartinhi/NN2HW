library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity RAM is
    port (
        in_ram_input_index: in std_logic_vector(7 downto 0); -- this is the given memory address
        out_data_ram:       out std_logic_vector(11 downto 0) -- this is the output datastream
    );
end RAM;

architecture RTL of RAM is
    type t_ram_arr is array (0 to 196) of std_logic_vector(11 downto 0);
    constant ram_arr: t_ram_arr := (
        -- here follows the generated array allocation
		"111000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110010000000",
		"000000011110",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"010000000000",
		"110110100110",
		"000011110110",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"011000000000",
		"100110110110",
		"011110110001",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110001000000",
		"000010110110",
		"100110100000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110100000000",
		"000010111110",
		"110101000000",
		"000000000010",
		"000000000000",
		"000000000000",
		"000000000000",
		"110100000000",
		"000001110110",
		"110100000000",
		"000000000101",
		"000000000000",
		"000000000000",
		"000000000000",
		"110100000000",
		"000000010110",
		"110010000000",
		"000000000110",
		"000000000000",
		"000000000000",
		"000000000000",
		"110110000000",
		"000000000110",
		"110001000000",
		"000000000110",
		"000000000000",
		"000000000000",
		"000000000000",
		"110110001000",
		"000000000110",
		"110001000000",
		"000000000110",
		"000000000000",
		"000000000000",
		"000000000000",
		"110110011000",
		"000000000110",
		"110001000000",
		"000000000110",
		"000000000000",
		"000000000000",
		"000000000000",
		"110110110000",
		"000000000100",
		"110001000000",
		"000000000110",
		"000000000000",
		"000000000000",
		"000000000000",
		"100110110000",
		"000000000000",
		"110001000000",
		"000000000110",
		"000000000000",
		"000000000000",
		"000000000000",
		"100110110000",
		"000000000000",
		"110011000000",
		"000000000101",
		"000000000000",
		"000000000000",
		"000000000000",
		"010110110000",
		"000000000000",
		"110100000000",
		"000000000001",
		"000000000000",
		"000000000000",
		"000000000000",
		"001110110000",
		"000000000000",
		"110101000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"100110110000",
		"000000000000",
		"100110100000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"100110100000",
		"001000000000",
		"000101110101",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110110000000",
		"110110100101",
		"000000101110",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"110011000000",
		"110110110110",
		"000000000101",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"001000000000",
		"010100110110",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000"

        -- here ends the generated array allocation
    );

begin
    out_data_ram <= ram_arr(to_integer(unsigned(in_ram_input_index)));
end RTL;

