library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
    port (
        reset:                  in std_logic;
        in_rom_input_index:     in std_logic_vector(7 downto 0); -- the given rom input index
        in_rom_neuron_index:    in std_logic_vector(3 downto 0); -- the given neuron index
        out_weights:            out std_logic_vector(31 downto 0) -- the output datastream
    );
end ROM;

architecture RTL of ROM is 
    type t_rom_arr is array (0 to 2500) of std_logic_vector (31 downto 0);
    signal rom_arr: t_rom_arr;

    signal rom_index: std_logic_vector (12 downto 0);
begin
    rom_index <= in_rom_neuron_index & in_rom_input_index; -- combine the neuron and input index to adress the array
    
    -- here follows the generated array allocation

    rom_arr(integer(2500)) <= "01110001011101010111100001111010";
    rom_arr(integer(2499)) <= "01110101011011010111011001110101";
    rom_arr(integer(2498)) <= "01111001011110000111011001110101";
    rom_arr(integer(2497)) <= "01110011011100010111100101110001";
    rom_arr(integer(2496)) <= "01110100011100100111011101110011";
    rom_arr(integer(2495)) <= "01110100011110010111010001111001";
    rom_arr(integer(2494)) <= "01110111011101010111100101110001";
    rom_arr(integer(2493)) <= "01110111011101000111100101111001";
    rom_arr(integer(2492)) <= "01110111011100010110110001101110";
    rom_arr(integer(2491)) <= "01110000011100010110110001101110";
    rom_arr(integer(2490)) <= "01101110011011100110101101110110";
    rom_arr(integer(2489)) <= "01110100011011100111000001101111";
    rom_arr(integer(2488)) <= "01110101011101100111011001110001";
    rom_arr(integer(2487)) <= "01110110011100010111011101110100";
    rom_arr(integer(2486)) <= "01110001011110000111100001111000";
    rom_arr(integer(2485)) <= "01110111011011010110011001100110";
    rom_arr(integer(2484)) <= "01100101010110110101101101100100";
    rom_arr(integer(2483)) <= "01011011010110110110000101011110";
    rom_arr(integer(2482)) <= "01100010010111010110011101100110";
    rom_arr(integer(2481)) <= "01101010011011000110111101110000";
    rom_arr(integer(2480)) <= "01110111011101000111011101111001";
    rom_arr(integer(2479)) <= "01110101011101100111001101110001";
    rom_arr(integer(2478)) <= "01110100011010000110010101011011";
    rom_arr(integer(2477)) <= "01100000011101001000001110000011";
    rom_arr(integer(2476)) <= "10001101100110001001101110011110";
    rom_arr(integer(2475)) <= "01110101100011001000011101111011";
    rom_arr(integer(2474)) <= "01101100011011100111001001110010";
    rom_arr(integer(2473)) <= "01110101011101000111100001110101";
    rom_arr(integer(2472)) <= "01110001011100100111010001101101";
    rom_arr(integer(2471)) <= "01101110011101000110100101100110";
    rom_arr(integer(2470)) <= "01101110011100001000111001110010";
    rom_arr(integer(2469)) <= "01111110100010011000011110000101";
    rom_arr(integer(2468)) <= "10011001100110011000111110000101";
    rom_arr(integer(2467)) <= "10001101011110000110100001100000";
    rom_arr(integer(2466)) <= "01110011011110010111011001110011";
    rom_arr(integer(2465)) <= "01110100011100010110111101101000";
    rom_arr(integer(2464)) <= "01110111100001000111011001111001";
    rom_arr(integer(2463)) <= "10000101011100111000101101111110";
    rom_arr(integer(2462)) <= "10000001011110011010100110000010";
    rom_arr(integer(2461)) <= "01110111100010101000100110001100";
    rom_arr(integer(2460)) <= "01111111100011001000000001011110";
    rom_arr(integer(2459)) <= "01110110011101010111011101110111";
    rom_arr(integer(2458)) <= "01110100011111010111001001101000";
    rom_arr(integer(2457)) <= "01101110011111110111101101111001";
    rom_arr(integer(2456)) <= "01110010011100110110111001111100";
    rom_arr(integer(2455)) <= "01111011011100000111010010010011";
    rom_arr(integer(2454)) <= "10001101100010100111110101111000";
    rom_arr(integer(2453)) <= "10010011100011001000011001110101";
    rom_arr(integer(2452)) <= "01110110011100010111011001110110";
    rom_arr(integer(2451)) <= "01110101011101000111001001101110";
    rom_arr(integer(2450)) <= "01101101100101011000100001111111";
    rom_arr(integer(2449)) <= "10000000011111101000000101101101";
    rom_arr(integer(2448)) <= "10000000011100101000100010100111";
    rom_arr(integer(2447)) <= "10010011100101111001001110010100";
    rom_arr(integer(2446)) <= "10001010100100001001010010000011";
    rom_arr(integer(2445)) <= "01101111011110010111010101110110";
    rom_arr(integer(2444)) <= "01111001011100110111000101110111";
    rom_arr(integer(2443)) <= "01111110100110011000110110000001";
    rom_arr(integer(2442)) <= "01101110100000110111111101101001";
    rom_arr(integer(2441)) <= "01101101011011000110100010011010";
    rom_arr(integer(2440)) <= "10011100100011010111101110010010";
    rom_arr(integer(2439)) <= "10010010100100111000001101111110";
    rom_arr(integer(2438)) <= "01101101011100010111011001110010";
    rom_arr(integer(2437)) <= "01110011011110000111000001111011";
    rom_arr(integer(2436)) <= "10000011100100100111010101101111";
    rom_arr(integer(2435)) <= "01110001011101010111101001110101";
    rom_arr(integer(2434)) <= "01110000011010000110000001101110";
    rom_arr(integer(2433)) <= "01111010101001111001011110011001";
    rom_arr(integer(2432)) <= "10000101100011000111111110000001";
    rom_arr(integer(2431)) <= "01110000011101010111100101111000";
    rom_arr(integer(2430)) <= "01110101011100010110111101111101";
    rom_arr(integer(2429)) <= "10000011100010110111100110001101";
    rom_arr(integer(2428)) <= "10000000011101001001110101110010";
    rom_arr(integer(2427)) <= "01101000011000100101111001110100";
    rom_arr(integer(2426)) <= "10000010101100001001011101111001";
    rom_arr(integer(2425)) <= "10001111100110011001000110000101";
    rom_arr(integer(2424)) <= "01110101011101000111100101110010";
    rom_arr(integer(2423)) <= "01110010011101000110101110000010";
    rom_arr(integer(2422)) <= "10001000100011001000100110010001";
    rom_arr(integer(2421)) <= "10000000100000101000001001101011";
    rom_arr(integer(2420)) <= "01101010010111000101100001101011";
    rom_arr(integer(2419)) <= "10010111100011001001000110011001";
    rom_arr(integer(2418)) <= "10001111100100001001010010001000";
    rom_arr(integer(2417)) <= "01110010011100110111100001110100";
    rom_arr(integer(2416)) <= "01110110011100000111110010011001";
    rom_arr(integer(2415)) <= "10010010100010001000001110010001";
    rom_arr(integer(2414)) <= "01110011011111100111000001100010";
    rom_arr(integer(2413)) <= "01011010010011100110010001110011";
    rom_arr(integer(2412)) <= "01101100100111111001000010010010";
    rom_arr(integer(2411)) <= "10011101011101001001100110001010";
    rom_arr(integer(2410)) <= "01100111011100000111100101110110";
    rom_arr(integer(2409)) <= "01111001011101111000010010100000";
    rom_arr(integer(2408)) <= "10011000100000111000111010000111";
    rom_arr(integer(2407)) <= "01110100011110000111000101011001";
    rom_arr(integer(2406)) <= "01011001010110000110110110101111";
    rom_arr(integer(2405)) <= "10011110011011101000111010000110";
    rom_arr(integer(2404)) <= "10100001100010001001001001110000";
    rom_arr(integer(2403)) <= "01101010011100100111011101110110";
    rom_arr(integer(2402)) <= "01110110011100011000000110011011";
    rom_arr(integer(2401)) <= "10010111100011010111110101101001";
    rom_arr(integer(2400)) <= "01111001011110010110111001011011";
    rom_arr(integer(2399)) <= "01010011010110010110011010000010";
    rom_arr(integer(2398)) <= "01111010100111010111111110001001";
    rom_arr(integer(2397)) <= "10010110100111010111100110000100";
    rom_arr(integer(2396)) <= "01110101011100110111101001110001";
    rom_arr(integer(2395)) <= "01111000011011100111000110101110";
    rom_arr(integer(2394)) <= "10010011100101001001000110010000";
    rom_arr(integer(2393)) <= "10001101011101000111001101011110";
    rom_arr(integer(2392)) <= "01011001011000011000011010101000";
    rom_arr(integer(2391)) <= "10000100100000110111111001111111";
    rom_arr(integer(2390)) <= "10001110101000010111011101110000";
    rom_arr(integer(2389)) <= "01110100011101000111010001111001";
    rom_arr(integer(2388)) <= "01110100011001110110011110010010";
    rom_arr(integer(2387)) <= "10001101100101001010000110001111";
    rom_arr(integer(2386)) <= "10000010011010010111001101011100";
    rom_arr(integer(2385)) <= "01011011011011001000001001101000";
    rom_arr(integer(2384)) <= "10001000011111110111001010001111";
    rom_arr(integer(2383)) <= "10010000100001110110111001101101";
    rom_arr(integer(2382)) <= "01110101011101100111001101111000";
    rom_arr(integer(2381)) <= "01110110011001010110000110100000";
    rom_arr(integer(2380)) <= "10011000100101001000100110001110";
    rom_arr(integer(2379)) <= "01110011100101101011011001111111";
    rom_arr(integer(2378)) <= "01101110100011111000110101111001";
    rom_arr(integer(2377)) <= "10001101011100111001001001111001";
    rom_arr(integer(2376)) <= "01111100011110011000011101110011";
    rom_arr(integer(2375)) <= "01111001011101110111000101110010";
    rom_arr(integer(2374)) <= "01110010011001110101111110100011";
    rom_arr(integer(2373)) <= "10011011011100110111011110001110";
    rom_arr(integer(2372)) <= "10011001100100111001000010001000";
    rom_arr(integer(2371)) <= "01100010011101011001111101110010";
    rom_arr(integer(2370)) <= "01110010100100100111110101110000";
    rom_arr(integer(2369)) <= "01110101011100010111011101110001";
    rom_arr(integer(2368)) <= "01111110011100100111100101110011";
    rom_arr(integer(2367)) <= "01110111011001100101011010001111";
    rom_arr(integer(2366)) <= "10101000100011001001000010010000";
    rom_arr(integer(2365)) <= "01110111100001111000111110101100";
    rom_arr(integer(2364)) <= "10001101100011100110111010001100";
    rom_arr(integer(2363)) <= "01110100011110101000111110000001";
    rom_arr(integer(2362)) <= "01111010011110100111010101101100";
    rom_arr(integer(2361)) <= "01110111011100010111010101111001";
    rom_arr(integer(2360)) <= "01110001011001000101110101110001";
    rom_arr(integer(2359)) <= "10010001011100110111110001111000";
    rom_arr(integer(2358)) <= "10001000100100101001010101110000";
    rom_arr(integer(2357)) <= "01110011011111001000011001110100";
    rom_arr(integer(2356)) <= "10001000100000101000100001110000";
    rom_arr(integer(2355)) <= "10000111100000110111011101110001";
    rom_arr(integer(2354)) <= "01110100011110000111001001110011";
    rom_arr(integer(2353)) <= "01110110011011000101110001011110";
    rom_arr(integer(2352)) <= "01110011100111111001100110001000";
    rom_arr(integer(2351)) <= "01111101100011101000000010001101";
    rom_arr(integer(2350)) <= "01110010100011111001000001101111";
    rom_arr(integer(2349)) <= "01110111011111000110100001111111";
    rom_arr(integer(2348)) <= "01111110100000010111000001101111";
    rom_arr(integer(2347)) <= "01111000011101110111001101110110";
    rom_arr(integer(2346)) <= "01110010011100000110011101100110";
    rom_arr(integer(2345)) <= "01101100011110101000000001110010";
    rom_arr(integer(2344)) <= "10001001100101011001001110000101";
    rom_arr(integer(2343)) <= "10000001100100001001000101110100";
    rom_arr(integer(2342)) <= "10010011100110011000010010000001";
    rom_arr(integer(2341)) <= "01111011011101010110010101110101";
    rom_arr(integer(2340)) <= "01110101011101100111011101110111";
    rom_arr(integer(2339)) <= "01111001011101000111000101101100";
    rom_arr(integer(2338)) <= "01110101011110100111010001111001";
    rom_arr(integer(2337)) <= "10000001100010111001011110000111";
    rom_arr(integer(2336)) <= "10011000100001011001011010001001";
    rom_arr(integer(2335)) <= "10100000011111111000011001111000";
    rom_arr(integer(2334)) <= "01110110011001110110101001110010";
    rom_arr(integer(2333)) <= "01110111011100010111100001110001";
    rom_arr(integer(2332)) <= "01110001011101000111011101110100";
    rom_arr(integer(2331)) <= "01110011011011010110100101110010";
    rom_arr(integer(2330)) <= "01110010011101101000101010001111";
    rom_arr(integer(2329)) <= "10000011100100011000111101111010";
    rom_arr(integer(2328)) <= "01111100011110110111010001110101";
    rom_arr(integer(2327)) <= "01100111011011010110111001111001";
    rom_arr(integer(2326)) <= "01111000011100100111011101110010";
    rom_arr(integer(2325)) <= "01110001011101010111010101111001";
    rom_arr(integer(2324)) <= "01110011011100100111000101101110";
    rom_arr(integer(2323)) <= "01110001011100000110110101101100";
    rom_arr(integer(2322)) <= "01100111011010110110111001110110";
    rom_arr(integer(2321)) <= "01110011011100100111010101110101";
    rom_arr(integer(2320)) <= "01110101011100010111100001111000";
    rom_arr(integer(2319)) <= "01111001011101010111100001110010";
    rom_arr(integer(2318)) <= "01110010011110010111010001110101";
    rom_arr(integer(2317)) <= "01110001011100010111011101110111";
    rom_arr(integer(2316)) <= "01111000011110010111101001111100";
    rom_arr(integer(2315)) <= "01110100011100000111100001111001";
    rom_arr(integer(2314)) <= "01110101011100010111011101111001";
    rom_arr(integer(2313)) <= "01110110011101100111001101110010";
    rom_arr(integer(2312)) <= "01111000011101110111010101110110";
    rom_arr(integer(2311)) <= "01110101011101100111100101110010";
    rom_arr(integer(2310)) <= "01111001011100010111010101110111";
    rom_arr(integer(2309)) <= "01110001011110010111100001110110";
    rom_arr(integer(2308)) <= "01110101011100110111011001110101";
    rom_arr(integer(2307)) <= "01110100011110000111001101110010";
    rom_arr(integer(2306)) <= "01111000011101010111011001110001";
    rom_arr(integer(2305)) <= "01110110011101000111001001111000";
    rom_arr(integer(2304)) <= "01010000000000000000000000000000";
    rom_arr(integer(2244)) <= "01110011011100010111010001110011";
    rom_arr(integer(2243)) <= "01110100011101110111011101110011";
    rom_arr(integer(2242)) <= "01110100011100000111000101110001";
    rom_arr(integer(2241)) <= "01111010011101110111000001110100";
    rom_arr(integer(2240)) <= "01111001011100010111100001110101";
    rom_arr(integer(2239)) <= "01110111011101100111001001110110";
    rom_arr(integer(2238)) <= "01110001011100010111010001110110";
    rom_arr(integer(2237)) <= "01110100011101100111011101110110";
    rom_arr(integer(2236)) <= "01110011011101000111001101110000";
    rom_arr(integer(2235)) <= "01101111011100000111001101101110";
    rom_arr(integer(2234)) <= "01110001011010010110100101101101";
    rom_arr(integer(2233)) <= "01101011011010110110111101101111";
    rom_arr(integer(2232)) <= "01110011011101100111001101110110";
    rom_arr(integer(2231)) <= "01110110011101000111100001110011";
    rom_arr(integer(2230)) <= "01110100011110010111011101111001";
    rom_arr(integer(2229)) <= "01111001011101000111100101101110";
    rom_arr(integer(2228)) <= "01101011011001100110000101011000";
    rom_arr(integer(2227)) <= "01100001011010000110110001101000";
    rom_arr(integer(2226)) <= "01011001010011010110101101101000";
    rom_arr(integer(2225)) <= "01101000011010110110011101110001";
    rom_arr(integer(2224)) <= "01110010011110000111100001110110";
    rom_arr(integer(2223)) <= "01110101011100100111100101110011";
    rom_arr(integer(2222)) <= "01110000011010110111010001110010";
    rom_arr(integer(2221)) <= "01111101011111010111100001010111";
    rom_arr(integer(2220)) <= "01110000011101000110011001101100";
    rom_arr(integer(2219)) <= "01100110011100010111100001101001";
    rom_arr(integer(2218)) <= "01110101011100110111010001101110";
    rom_arr(integer(2217)) <= "01110000011100110111001001110010";
    rom_arr(integer(2216)) <= "01110111011110110111010001110101";
    rom_arr(integer(2215)) <= "01101011011011100110011001111010";
    rom_arr(integer(2214)) <= "10000110011100101001100101111110";
    rom_arr(integer(2213)) <= "10000101011010001000001110010010";
    rom_arr(integer(2212)) <= "10000011011110001000010001111111";
    rom_arr(integer(2211)) <= "10000010100011011000110001101100";
    rom_arr(integer(2210)) <= "01101010011101110111101001110111";
    rom_arr(integer(2209)) <= "01110010011101110111011001111011";
    rom_arr(integer(2208)) <= "01110000011001011000010110011111";
    rom_arr(integer(2207)) <= "10011000101001101001010101111011";
    rom_arr(integer(2206)) <= "01111010011101110101001000111111";
    rom_arr(integer(2205)) <= "01011111011101001000010110000110";
    rom_arr(integer(2204)) <= "10001000101001101100011010000101";
    rom_arr(integer(2203)) <= "01111010011101010111001001110100";
    rom_arr(integer(2202)) <= "01111001011110010111100110001000";
    rom_arr(integer(2201)) <= "01101110011001111001011010100010";
    rom_arr(integer(2200)) <= "10001101101001010110111001110101";
    rom_arr(integer(2199)) <= "10001010100010010111110110000000";
    rom_arr(integer(2198)) <= "01111111100100001000010010001010";
    rom_arr(integer(2197)) <= "10011011101000001010001110000001";
    rom_arr(integer(2196)) <= "01111111011100100111010001110101";
    rom_arr(integer(2195)) <= "01111001011110110111110010000000";
    rom_arr(integer(2194)) <= "01110101011110101000110110010010";
    rom_arr(integer(2193)) <= "10011100101011001010011110011000";
    rom_arr(integer(2192)) <= "01101110011110000111010110000011";
    rom_arr(integer(2191)) <= "10001100100100001000101110010111";
    rom_arr(integer(2190)) <= "10001100011110000101001101110000";
    rom_arr(integer(2189)) <= "01110111011101110111100001110100";
    rom_arr(integer(2188)) <= "01110100011110010111110110001010";
    rom_arr(integer(2187)) <= "01111111011110000111010110001000";
    rom_arr(integer(2186)) <= "10010110011111100110100110011001";
    rom_arr(integer(2185)) <= "10000000011101011000011001111000";
    rom_arr(integer(2184)) <= "01111001100001111001000101111011";
    rom_arr(integer(2183)) <= "10001000011011000101001001101001";
    rom_arr(integer(2182)) <= "01110100011101010111010001110100";
    rom_arr(integer(2181)) <= "01110011011101100111101010000001";
    rom_arr(integer(2180)) <= "01111001011110001000001110001110";
    rom_arr(integer(2179)) <= "01110100011110000111000101011000";
    rom_arr(integer(2178)) <= "01100011100100011000110010000100";
    rom_arr(integer(2177)) <= "01110101011110001000010010000101";
    rom_arr(integer(2176)) <= "01101000010100010101110101110100";
    rom_arr(integer(2175)) <= "01111000011101100111010001110101";
    rom_arr(integer(2174)) <= "01111001011100100111000001111010";
    rom_arr(integer(2173)) <= "01110111011111010111010001110100";
    rom_arr(integer(2172)) <= "01101110011010110101101001100110";
    rom_arr(integer(2171)) <= "10000010100101101001000110001001";
    rom_arr(integer(2170)) <= "01110011100010110111010101110110";
    rom_arr(integer(2169)) <= "01101011010111100110011101110001";
    rom_arr(integer(2168)) <= "01110000011101010111000001111001";
    rom_arr(integer(2167)) <= "01110110011101100111000001111001";
    rom_arr(integer(2166)) <= "01101011011010100111001101101001";
    rom_arr(integer(2165)) <= "01011101010111010101011101111010";
    rom_arr(integer(2164)) <= "01110000101010011001001001110110";
    rom_arr(integer(2163)) <= "01111010011101101000010101110101";
    rom_arr(integer(2162)) <= "01101011011001100111000101111000";
    rom_arr(integer(2161)) <= "01110101011110100111100001110101";
    rom_arr(integer(2160)) <= "01110011011101110111011101110001";
    rom_arr(integer(2159)) <= "01101111011011100111000001011111";
    rom_arr(integer(2158)) <= "01010110010111100110011010100011";
    rom_arr(integer(2157)) <= "10000101101011001001010010010010";
    rom_arr(integer(2156)) <= "01111000011010000110111010000101";
    rom_arr(integer(2155)) <= "01110010011010100110110101110111";
    rom_arr(integer(2154)) <= "01110010011110010111100001110010";
    rom_arr(integer(2153)) <= "01110101011110010110111101110010";
    rom_arr(integer(2152)) <= "01101111011011110110111001101100";
    rom_arr(integer(2151)) <= "01011111011000110110111110000101";
    rom_arr(integer(2150)) <= "10010010101000111001000110001000";
    rom_arr(integer(2149)) <= "01100101010110110111000010000001";
    rom_arr(integer(2148)) <= "01101010011100110111010001110111";
    rom_arr(integer(2147)) <= "01111001011100110111000101111001";
    rom_arr(integer(2146)) <= "01110110011101010111001001101100";
    rom_arr(integer(2145)) <= "01110000011011110111010101101111";
    rom_arr(integer(2144)) <= "01101000011011101010000010000111";
    rom_arr(integer(2143)) <= "10010101101000101001010110001011";
    rom_arr(integer(2142)) <= "01100111010110110111100110001000";
    rom_arr(integer(2141)) <= "01110111011101100111100101111100";
    rom_arr(integer(2140)) <= "01110101011110000111011001111000";
    rom_arr(integer(2139)) <= "01110111011101010111010101110000";
    rom_arr(integer(2138)) <= "01110110011101110111011101110101";
    rom_arr(integer(2137)) <= "01101110011101101000000110001010";
    rom_arr(integer(2136)) <= "10011110101011011001100010000111";
    rom_arr(integer(2135)) <= "01101111011100100111110101110101";
    rom_arr(integer(2134)) <= "01111100011110000111010001110101";
    rom_arr(integer(2133)) <= "01111000011100010111100001110001";
    rom_arr(integer(2132)) <= "01110010011101100111001101100110";
    rom_arr(integer(2131)) <= "01101100011010010111000101110110";
    rom_arr(integer(2130)) <= "01110101011111100111001110010000";
    rom_arr(integer(2129)) <= "10101011101010001001110101111010";
    rom_arr(integer(2128)) <= "01110101011101110111001101110010";
    rom_arr(integer(2127)) <= "01101010010110100110101101110000";
    rom_arr(integer(2126)) <= "01110100011101110111011001110110";
    rom_arr(integer(2125)) <= "01111001011101110110110101100011";
    rom_arr(integer(2124)) <= "01100001011001110111011101101010";
    rom_arr(integer(2123)) <= "01110111011100111000100010010001";
    rom_arr(integer(2122)) <= "10101000100100111001001001111001";
    rom_arr(integer(2121)) <= "10001101011110110111001001111000";
    rom_arr(integer(2120)) <= "01101000010110010101101001100111";
    rom_arr(integer(2119)) <= "01110100011101100111100101110010";
    rom_arr(integer(2118)) <= "01111000011100010110011101100101";
    rom_arr(integer(2117)) <= "01100010011011010111001101101011";
    rom_arr(integer(2116)) <= "01101110011110011000000110001101";
    rom_arr(integer(2115)) <= "10010010100010000111101101110001";
    rom_arr(integer(2114)) <= "01110011011100110111000001110100";
    rom_arr(integer(2113)) <= "01110101011001010101100001101101";
    rom_arr(integer(2112)) <= "01111000011101100111011001111001";
    rom_arr(integer(2111)) <= "01111001011011110110011001010010";
    rom_arr(integer(2110)) <= "01011111011100010110111001101100";
    rom_arr(integer(2109)) <= "01111101011101101000011001101010";
    rom_arr(integer(2108)) <= "10000100011111000111110001111001";
    rom_arr(integer(2107)) <= "01101010011100010110011101101000";
    rom_arr(integer(2106)) <= "01101111011000100110010101110110";
    rom_arr(integer(2105)) <= "01111000011011010111001001110011";
    rom_arr(integer(2104)) <= "01110010011101100110001001011100";
    rom_arr(integer(2103)) <= "01110001011101101000000010000100";
    rom_arr(integer(2102)) <= "01111111011100000110111001111000";
    rom_arr(integer(2101)) <= "01011000011111000110100110000000";
    rom_arr(integer(2100)) <= "01101101011100100110111101100001";
    rom_arr(integer(2099)) <= "01101111011000000110011001111001";
    rom_arr(integer(2098)) <= "01110100011011110111000101110101";
    rom_arr(integer(2097)) <= "01110101011101110110010101111001";
    rom_arr(integer(2096)) <= "10000001011111100111110101111111";
    rom_arr(integer(2095)) <= "01101010100000000101101001110011";
    rom_arr(integer(2094)) <= "01100001011010100110110101110000";
    rom_arr(integer(2093)) <= "01110111011100100110101001101000";
    rom_arr(integer(2092)) <= "01100111011100010111010101110110";
    rom_arr(integer(2091)) <= "01110011011100000111011101110101";
    rom_arr(integer(2090)) <= "01110111011011110110001101101110";
    rom_arr(integer(2089)) <= "01111111100010101000100001111111";
    rom_arr(integer(2088)) <= "01111101011111010110101001111100";
    rom_arr(integer(2087)) <= "10000101011101010111101001101101";
    rom_arr(integer(2086)) <= "01101010011100010110100001100111";
    rom_arr(integer(2085)) <= "01111001100001001000000001111010";
    rom_arr(integer(2084)) <= "01111010011110000111001001110111";
    rom_arr(integer(2083)) <= "01110110011100110110100101010101";
    rom_arr(integer(2082)) <= "01101010011011010111100101111110";
    rom_arr(integer(2081)) <= "10000011011111001000001110001010";
    rom_arr(integer(2080)) <= "10000111100010101001000110000011";
    rom_arr(integer(2079)) <= "01110110011110010111001101111100";
    rom_arr(integer(2078)) <= "01110010011111100111101001110001";
    rom_arr(integer(2077)) <= "01110010011101110111100001110100";
    rom_arr(integer(2076)) <= "01110011011101010111011101110000";
    rom_arr(integer(2075)) <= "01101111011011010110101001110010";
    rom_arr(integer(2074)) <= "01110100011001110111011010001101";
    rom_arr(integer(2073)) <= "10000100011101000111110001110101";
    rom_arr(integer(2072)) <= "01100010011001100110111001110000";
    rom_arr(integer(2071)) <= "01110100011101000111100001110100";
    rom_arr(integer(2070)) <= "01110111011100000111011001110011";
    rom_arr(integer(2069)) <= "01111001011110000111100101110101";
    rom_arr(integer(2068)) <= "01111001011100110111000101111000";
    rom_arr(integer(2067)) <= "01110100011110000111011010001000";
    rom_arr(integer(2066)) <= "10010010011111111000001101110001";
    rom_arr(integer(2065)) <= "01110000011011010110111101110101";
    rom_arr(integer(2064)) <= "01110100011100100111100001110100";
    rom_arr(integer(2063)) <= "01110110011101100111100101111000";
    rom_arr(integer(2062)) <= "01111001011100100111001101110001";
    rom_arr(integer(2061)) <= "01110101011101000111000101111001";
    rom_arr(integer(2060)) <= "01111010011101010111001101110100";
    rom_arr(integer(2059)) <= "01111010011110100111011101110001";
    rom_arr(integer(2058)) <= "01111010011110000111011001110100";
    rom_arr(integer(2057)) <= "01110010011101110111010101111000";
    rom_arr(integer(2056)) <= "01110111011101000111100001110011";
    rom_arr(integer(2055)) <= "01110110011110010111010001110111";
    rom_arr(integer(2054)) <= "01110100011100010111011101110111";
    rom_arr(integer(2053)) <= "01111000011101110111000101110111";
    rom_arr(integer(2052)) <= "01111000011101110111000101110001";
    rom_arr(integer(2051)) <= "01110110011100010111000101110100";
    rom_arr(integer(2050)) <= "01110010011110010111001001110011";
    rom_arr(integer(2049)) <= "01111000011101000111010001110111";
    rom_arr(integer(2048)) <= "10111001000000000000000000000000";
    rom_arr(integer(1988)) <= "01110101011100010111100001110110";
    rom_arr(integer(1987)) <= "01110110011101100111011001110110";
    rom_arr(integer(1986)) <= "01110111011101100111010001110010";
    rom_arr(integer(1985)) <= "01110110011101000111100101111000";
    rom_arr(integer(1984)) <= "01111010011100010111011101110110";
    rom_arr(integer(1983)) <= "01110100011110000111100101111000";
    rom_arr(integer(1982)) <= "01110001011101010111010001110100";
    rom_arr(integer(1981)) <= "01111000011100010111010101110001";
    rom_arr(integer(1980)) <= "01110101011100110111001101110100";
    rom_arr(integer(1979)) <= "01110010011011010110110001101110";
    rom_arr(integer(1978)) <= "01101100011011100110111001110000";
    rom_arr(integer(1977)) <= "01110001011101000111011101101110";
    rom_arr(integer(1976)) <= "01110000011110010111000001110110";
    rom_arr(integer(1975)) <= "01111000011110000111001101110111";
    rom_arr(integer(1974)) <= "01111000011111000111011001111000";
    rom_arr(integer(1973)) <= "01110010011001010110010101100100";
    rom_arr(integer(1972)) <= "01100101011011100111111110001000";
    rom_arr(integer(1971)) <= "10010101100010110111010101110100";
    rom_arr(integer(1970)) <= "01101000011001110101110001011110";
    rom_arr(integer(1969)) <= "01101010011011110110111001110001";
    rom_arr(integer(1968)) <= "01101111011101000111011101110100";
    rom_arr(integer(1967)) <= "01110011011110001000100110010111";
    rom_arr(integer(1966)) <= "10000000100000001000111010000000";
    rom_arr(integer(1965)) <= "10000100101001101010101001110010";
    rom_arr(integer(1964)) <= "01101011111111110110010010100000";
    rom_arr(integer(1963)) <= "01110111011111111000101101111001";
    rom_arr(integer(1962)) <= "01101111011001110110000101101101";
    rom_arr(integer(1961)) <= "01101010011100100111010101110111";
    rom_arr(integer(1960)) <= "01110110011101010111111110001100";
    rom_arr(integer(1959)) <= "10010001100111001001111110010001";
    rom_arr(integer(1958)) <= "10101011101001010110111110001001";
    rom_arr(integer(1957)) <= "01101110011100100110101010001101";
    rom_arr(integer(1956)) <= "10010010011011111001011101111001";
    rom_arr(integer(1955)) <= "10010011011111110111011001111001";
    rom_arr(integer(1954)) <= "01110110011110010111000101110010";
    rom_arr(integer(1953)) <= "01110011011100011000000010000110";
    rom_arr(integer(1952)) <= "10000011100011001000000010010100";
    rom_arr(integer(1951)) <= "01111000100011010111000101111110";
    rom_arr(integer(1950)) <= "01110010011110000111101001111011";
    rom_arr(integer(1949)) <= "01111111100000001001101110100011";
    rom_arr(integer(1948)) <= "10100011100111111000010110001110";
    rom_arr(integer(1947)) <= "10000010011111110111011101110110";
    rom_arr(integer(1946)) <= "01110101011101111000011010000111";
    rom_arr(integer(1945)) <= "10011111100100111000110001111101";
    rom_arr(integer(1944)) <= "10111100100011011010010010000111";
    rom_arr(integer(1943)) <= "01101100011111111000101001110001";
    rom_arr(integer(1942)) <= "10000111100000011001100001100110";
    rom_arr(integer(1941)) <= "10000101100010111000000110000011";
    rom_arr(integer(1940)) <= "10000010100000110111100001110101";
    rom_arr(integer(1939)) <= "01110100011110011000011110010100";
    rom_arr(integer(1938)) <= "10001000100011111001110110100000";
    rom_arr(integer(1937)) <= "10011000100001100110110101111010";
    rom_arr(integer(1936)) <= "10000101011011100111101010000110";
    rom_arr(integer(1935)) <= "10101100100010101001110110010111";
    rom_arr(integer(1934)) <= "10111100100111101001011110010010";
    rom_arr(integer(1933)) <= "10000001100000000111001001110111";
    rom_arr(integer(1932)) <= "01111010100001001010100110000100";
    rom_arr(integer(1931)) <= "10001111100111111000110110000010";
    rom_arr(integer(1930)) <= "01101100100010011000111110001100";
    rom_arr(integer(1929)) <= "10001010011111011010011101111100";
    rom_arr(integer(1928)) <= "10000000101000001001101010001011";
    rom_arr(integer(1927)) <= "10001100011110001000101010001111";
    rom_arr(integer(1926)) <= "01101100011100100111011101110100";
    rom_arr(integer(1925)) <= "01110111011110101010100010101111";
    rom_arr(integer(1924)) <= "10100001100100101000100101110100";
    rom_arr(integer(1923)) <= "10001110011110011001101110000000";
    rom_arr(integer(1922)) <= "01101111100001011000001010110110";
    rom_arr(integer(1921)) <= "10000000100100110111100101111111";
    rom_arr(integer(1920)) <= "10101100100101111010111110010101";
    rom_arr(integer(1919)) <= "10000000011101110111001001110001";
    rom_arr(integer(1918)) <= "01111101100100111100100110001101";
    rom_arr(integer(1917)) <= "01110000011111110111010101111011";
    rom_arr(integer(1916)) <= "01111011011111100110011001110101";
    rom_arr(integer(1915)) <= "10010010011110011000110110001101";
    rom_arr(integer(1914)) <= "10001100101100011000110101111111";
    rom_arr(integer(1913)) <= "10010010100101001000101010010011";
    rom_arr(integer(1912)) <= "10010011100000000111001101110100";
    rom_arr(integer(1911)) <= "01111101101011111100000010100000";
    rom_arr(integer(1910)) <= "10001111101000001011101101101101";
    rom_arr(integer(1909)) <= "10001010011101001100011101111101";
    rom_arr(integer(1908)) <= "01110011100011101010000110010110";
    rom_arr(integer(1907)) <= "10001011100000001001111001101110";
    rom_arr(integer(1906)) <= "01111111100111101000010010011101";
    rom_arr(integer(1905)) <= "10011001011100110111001001111000";
    rom_arr(integer(1904)) <= "10000000100110111010011010100101";
    rom_arr(integer(1903)) <= "01101001011001110110111101101100";
    rom_arr(integer(1902)) <= "10000000011011110110101001111100";
    rom_arr(integer(1901)) <= "10000101011111101000011101111000";
    rom_arr(integer(1900)) <= "10001000011111011000000110001100";
    rom_arr(integer(1899)) <= "01111100101000011010000010001001";
    rom_arr(integer(1898)) <= "01110111011100010111011001110101";
    rom_arr(integer(1897)) <= "01111001100110001001110010010000";
    rom_arr(integer(1896)) <= "10001101011100110110111110001111";
    rom_arr(integer(1895)) <= "01110100100011010110101101111110";
    rom_arr(integer(1894)) <= "01110111100000011001000001111100";
    rom_arr(integer(1893)) <= "10001101100000100110111101110000";
    rom_arr(integer(1892)) <= "10000100011010000101010001010111";
    rom_arr(integer(1891)) <= "01101000011101010111100001110011";
    rom_arr(integer(1890)) <= "10001001101010001011000110111001";
    rom_arr(integer(1889)) <= "01111001100000011000111001101111";
    rom_arr(integer(1888)) <= "01101111011010010111011101110110";
    rom_arr(integer(1887)) <= "01101001011111001010001001111010";
    rom_arr(integer(1886)) <= "10010010011011010110101101101101";
    rom_arr(integer(1885)) <= "01011100010011010100001101000101";
    rom_arr(integer(1884)) <= "01100101011110010111011101110011";
    rom_arr(integer(1883)) <= "01110111100011101010001010000101";
    rom_arr(integer(1882)) <= "01100111011110111000111101111110";
    rom_arr(integer(1881)) <= "10010101011001010110101001110010";
    rom_arr(integer(1880)) <= "01100110011001100110100001101000";
    rom_arr(integer(1879)) <= "01100011011010000110100101101010";
    rom_arr(integer(1878)) <= "01011010010101000110010001100101";
    rom_arr(integer(1877)) <= "01100110011101100111001101111001";
    rom_arr(integer(1876)) <= "01110100011110000111110101101110";
    rom_arr(integer(1875)) <= "01110100011111101000101101110100";
    rom_arr(integer(1874)) <= "10011100011100110110001101110011";
    rom_arr(integer(1873)) <= "01101000011001000101110101100001";
    rom_arr(integer(1872)) <= "01100011010111010110101001101100";
    rom_arr(integer(1871)) <= "01110101100000001000000001101111";
    rom_arr(integer(1870)) <= "01110010011101110111010101110111";
    rom_arr(integer(1869)) <= "01111000011110100111000101011010";
    rom_arr(integer(1868)) <= "01110100011101001000000110000110";
    rom_arr(integer(1867)) <= "01110011100000001001101101111011";
    rom_arr(integer(1866)) <= "01101000011100100110110001111101";
    rom_arr(integer(1865)) <= "10000000011101010110111101111110";
    rom_arr(integer(1864)) <= "01111110101100111001101101101101";
    rom_arr(integer(1863)) <= "01111011011011110111011101111001";
    rom_arr(integer(1862)) <= "01110110011100010110100101011010";
    rom_arr(integer(1861)) <= "01111110100010110111010101111011";
    rom_arr(integer(1860)) <= "01110110100011000111101110001110";
    rom_arr(integer(1859)) <= "10010110100011110111011001111010";
    rom_arr(integer(1858)) <= "01101100100010011001010001110010";
    rom_arr(integer(1857)) <= "01110010011001011001111110001001";
    rom_arr(integer(1856)) <= "01111000011101100111000001110100";
    rom_arr(integer(1855)) <= "01110101011100100110011101011011";
    rom_arr(integer(1854)) <= "10000001011111010111001110001001";
    rom_arr(integer(1853)) <= "10100001011001111000011101110011";
    rom_arr(integer(1852)) <= "01111000011101100111000001101110";
    rom_arr(integer(1851)) <= "10000000100110110110111010000011";
    rom_arr(integer(1850)) <= "10000111011110011000000110010111";
    rom_arr(integer(1849)) <= "01111001011100110111010101110100";
    rom_arr(integer(1848)) <= "01110101011100010111001001011110";
    rom_arr(integer(1847)) <= "01011001100111011000000001101100";
    rom_arr(integer(1846)) <= "01101100011111010110010001111110";
    rom_arr(integer(1845)) <= "01101110011110111001101101101110";
    rom_arr(integer(1844)) <= "10000110011011100111010110011100";
    rom_arr(integer(1843)) <= "01110010100100011000100010011001";
    rom_arr(integer(1842)) <= "01111001011111000111011001110111";
    rom_arr(integer(1841)) <= "01110011011100010111001101100000";
    rom_arr(integer(1840)) <= "01011111011011100111001001110000";
    rom_arr(integer(1839)) <= "01110100011111010111010010000100";
    rom_arr(integer(1838)) <= "10000000011101100111110101111100";
    rom_arr(integer(1837)) <= "01110001100110011001010101110111";
    rom_arr(integer(1836)) <= "10001000011111010111101110000010";
    rom_arr(integer(1835)) <= "01110111011100100111001101110110";
    rom_arr(integer(1834)) <= "01110011011101110111001101100011";
    rom_arr(integer(1833)) <= "01101100011101100111111110001101";
    rom_arr(integer(1832)) <= "10000011100000101000010110011010";
    rom_arr(integer(1831)) <= "01111110100000001000100010001111";
    rom_arr(integer(1830)) <= "10011100011111100111101010001100";
    rom_arr(integer(1829)) <= "01111111011110000111110001110011";
    rom_arr(integer(1828)) <= "01110111011101110111100101110100";
    rom_arr(integer(1827)) <= "01110111011100010111011001100110";
    rom_arr(integer(1826)) <= "01011111011000000110110001110111";
    rom_arr(integer(1825)) <= "01111101100100101001101110100000";
    rom_arr(integer(1824)) <= "10010101101110001001000010101000";
    rom_arr(integer(1823)) <= "10100110100110001001101010000110";
    rom_arr(integer(1822)) <= "10000110100011110111010001101111";
    rom_arr(integer(1821)) <= "01110110011101100111010101110111";
    rom_arr(integer(1820)) <= "01110101011110000111001101110010";
    rom_arr(integer(1819)) <= "01101101011011100110111101101110";
    rom_arr(integer(1818)) <= "01110100011100111000100110010110";
    rom_arr(integer(1817)) <= "10000111100100001010001110001111";
    rom_arr(integer(1816)) <= "10010111100101011001110010000000";
    rom_arr(integer(1815)) <= "01111101011100100111100001111001";
    rom_arr(integer(1814)) <= "01110110011100100111000101110010";
    rom_arr(integer(1813)) <= "01111001011100100111100101111010";
    rom_arr(integer(1812)) <= "01110000011101000111010001110010";
    rom_arr(integer(1811)) <= "01101111011100101000000001111101";
    rom_arr(integer(1810)) <= "10001010011101110111101010000110";
    rom_arr(integer(1809)) <= "10000011011111111000001101110100";
    rom_arr(integer(1808)) <= "01110011011100110111011001110100";
    rom_arr(integer(1807)) <= "01110010011101110111001001110101";
    rom_arr(integer(1806)) <= "01110001011100110111010001110111";
    rom_arr(integer(1805)) <= "01110100011110000111001101110010";
    rom_arr(integer(1804)) <= "01111000011100110111001110000010";
    rom_arr(integer(1803)) <= "01111110011101100111001001101111";
    rom_arr(integer(1802)) <= "01110111011011110111011101110011";
    rom_arr(integer(1801)) <= "01110111011101100111100001110111";
    rom_arr(integer(1800)) <= "01110100011100100111011101111001";
    rom_arr(integer(1799)) <= "01111010011101010111000101111001";
    rom_arr(integer(1798)) <= "01111000011110000111101001110010";
    rom_arr(integer(1797)) <= "01111010011101110111001101110110";
    rom_arr(integer(1796)) <= "01111001011100100111001001111000";
    rom_arr(integer(1795)) <= "01110100011100010111010101110100";
    rom_arr(integer(1794)) <= "01111001011110000111100101111010";
    rom_arr(integer(1793)) <= "01110110011100100111001001110111";
    rom_arr(integer(1792)) <= "10000011000000000000000000000000";
    rom_arr(integer(1732)) <= "01110001011110010111001001110110";
    rom_arr(integer(1731)) <= "01110100011101010111101001110100";
    rom_arr(integer(1730)) <= "01110110011100100111010101110011";
    rom_arr(integer(1729)) <= "01111000011100100111000101110111";
    rom_arr(integer(1728)) <= "01110101011101000111001001110111";
    rom_arr(integer(1727)) <= "01110010011110000111100101110101";
    rom_arr(integer(1726)) <= "01111000011101100111100101111001";
    rom_arr(integer(1725)) <= "01111010011100010111000101110101";
    rom_arr(integer(1724)) <= "01111001011110010111001101111001";
    rom_arr(integer(1723)) <= "01111011100001101000100110010000";
    rom_arr(integer(1722)) <= "01111110100001001000110101111100";
    rom_arr(integer(1721)) <= "10001010011111100111010001111000";
    rom_arr(integer(1720)) <= "01110111011110010111011001110000";
    rom_arr(integer(1719)) <= "01111000011100010111011101111000";
    rom_arr(integer(1718)) <= "01110111011100010111011101110101";
    rom_arr(integer(1717)) <= "01110001011101110111001001111010";
    rom_arr(integer(1716)) <= "10100010100111001001110110101101";
    rom_arr(integer(1715)) <= "10100011100011111100100111010011";
    rom_arr(integer(1714)) <= "10101100101111001100000111001011";
    rom_arr(integer(1713)) <= "10100110100110011000000101111000";
    rom_arr(integer(1712)) <= "01101011011110100111010001111001";
    rom_arr(integer(1711)) <= "01110010011100010111001001110000";
    rom_arr(integer(1710)) <= "01110011011110001000000101111100";
    rom_arr(integer(1709)) <= "01110011011011011010000010100101";
    rom_arr(integer(1708)) <= "01111101101100011001110010000000";
    rom_arr(integer(1707)) <= "10011111100111100111111110001011";
    rom_arr(integer(1706)) <= "10011110101000101000010010011000";
    rom_arr(integer(1705)) <= "10001010011110010111100101110001";
    rom_arr(integer(1704)) <= "01111000011101010111001001101111";
    rom_arr(integer(1703)) <= "01101101011011100111010010000100";
    rom_arr(integer(1702)) <= "01111111101110010111001001101000";
    rom_arr(integer(1701)) <= "01111000011011011001000101101000";
    rom_arr(integer(1700)) <= "10010110100010111000101110000000";
    rom_arr(integer(1699)) <= "10010101100011111000110010011010";
    rom_arr(integer(1698)) <= "10010100100000010111011001110011";
    rom_arr(integer(1697)) <= "01111010011101000110111101101101";
    rom_arr(integer(1696)) <= "01110000100001110111010110011000";
    rom_arr(integer(1695)) <= "01111111011101011001010001111110";
    rom_arr(integer(1694)) <= "10001000011011100110111101101111";
    rom_arr(integer(1693)) <= "10001010011101111000001101111101";
    rom_arr(integer(1692)) <= "10001101100011000111100110000110";
    rom_arr(integer(1691)) <= "10001011011111110111010101111000";
    rom_arr(integer(1690)) <= "01110000011100100111011001100110";
    rom_arr(integer(1689)) <= "01110010100000100111000101101101";
    rom_arr(integer(1688)) <= "10101100100011110111101110000111";
    rom_arr(integer(1687)) <= "01111101011100010111010101110101";
    rom_arr(integer(1686)) <= "01110101011101100110011110001011";
    rom_arr(integer(1685)) <= "10011001100100010111000010001101";
    rom_arr(integer(1684)) <= "10001110011110000111011101110100";
    rom_arr(integer(1683)) <= "01110001011101000110111101110010";
    rom_arr(integer(1682)) <= "10001110100000011001001110111110";
    rom_arr(integer(1681)) <= "01111011100110111000101001111110";
    rom_arr(integer(1680)) <= "01110101100001100111001101100011";
    rom_arr(integer(1679)) <= "01111001011111111010110110001111";
    rom_arr(integer(1678)) <= "10010011101011101001100010011001";
    rom_arr(integer(1677)) <= "10010110011100100111001101111001";
    rom_arr(integer(1676)) <= "01110110011100110110110101110010";
    rom_arr(integer(1675)) <= "10011000011110011000110001110010";
    rom_arr(integer(1674)) <= "10001111100010101001011101111110";
    rom_arr(integer(1673)) <= "01110101011110010111110001110011";
    rom_arr(integer(1672)) <= "01110000100000110111010110000001";
    rom_arr(integer(1671)) <= "01110101011101111010000010001101";
    rom_arr(integer(1670)) <= "10010111011011010111000001111001";
    rom_arr(integer(1669)) <= "01110011011101110110110001100110";
    rom_arr(integer(1668)) <= "01111111101001101001111101111110";
    rom_arr(integer(1667)) <= "10000000011111111000001010100000";
    rom_arr(integer(1666)) <= "10001001011001110110101101101000";
    rom_arr(integer(1665)) <= "01101111011011010110100101111010";
    rom_arr(integer(1664)) <= "01111000101010001001100010001110";
    rom_arr(integer(1663)) <= "10100100011110010111001101110010";
    rom_arr(integer(1662)) <= "01110011011011110110010101101110";
    rom_arr(integer(1661)) <= "10011110100001010111111001110010";
    rom_arr(integer(1660)) <= "10100000011101101001100101110110";
    rom_arr(integer(1659)) <= "01100101011001000110011001100111";
    rom_arr(integer(1658)) <= "01101001011010000110011101110001";
    rom_arr(integer(1657)) <= "10001010011101011000010110100001";
    rom_arr(integer(1656)) <= "10010010011110100111100101110100";
    rom_arr(integer(1655)) <= "01110011011100100110100110100111";
    rom_arr(integer(1654)) <= "10100111100101101000000010001100";
    rom_arr(integer(1653)) <= "10010010100110000111110001100110";
    rom_arr(integer(1652)) <= "01110100011101001011111101110001";
    rom_arr(integer(1651)) <= "01111111011110110111101001100111";
    rom_arr(integer(1650)) <= "01101111011100101001000010010101";
    rom_arr(integer(1649)) <= "01111111011111110111010001111000";
    rom_arr(integer(1648)) <= "01110110011100100110111010010000";
    rom_arr(integer(1647)) <= "10100010100100101001000010100111";
    rom_arr(integer(1646)) <= "01111100011011100111111001111111";
    rom_arr(integer(1645)) <= "10001100100001110111001010000110";
    rom_arr(integer(1644)) <= "10000000011100100110111101101000";
    rom_arr(integer(1643)) <= "01101110011110000111000001111001";
    rom_arr(integer(1642)) <= "01111000011101010111100101110001";
    rom_arr(integer(1641)) <= "01110100011100010110111101110110";
    rom_arr(integer(1640)) <= "01110010011010010111111001101111";
    rom_arr(integer(1639)) <= "01101000100000100111111001111100";
    rom_arr(integer(1638)) <= "10000001100001011000010010010101";
    rom_arr(integer(1637)) <= "01110011011110110111101001110100";
    rom_arr(integer(1636)) <= "01101111011010110110011001101011";
    rom_arr(integer(1635)) <= "01111100011110010111011001110110";
    rom_arr(integer(1634)) <= "01110010011110010111101101110000";
    rom_arr(integer(1633)) <= "01100111010101010110100101110001";
    rom_arr(integer(1632)) <= "01111100100010110111101110001010";
    rom_arr(integer(1631)) <= "01110000100100001001111010001100";
    rom_arr(integer(1630)) <= "01111011011100100111001001110011";
    rom_arr(integer(1629)) <= "01110110011101000110111101101000";
    rom_arr(integer(1628)) <= "01110111011110010111010001110100";
    rom_arr(integer(1627)) <= "01110001011100010111100001101100";
    rom_arr(integer(1626)) <= "01100101011010000110100101111010";
    rom_arr(integer(1625)) <= "01110111100001110111011010001110";
    rom_arr(integer(1624)) <= "10000110100111110111111010010100";
    rom_arr(integer(1623)) <= "01111000101000000111001101101111";
    rom_arr(integer(1622)) <= "01111000011100010111000101110110";
    rom_arr(integer(1621)) <= "10000000011100000111000101110111";
    rom_arr(integer(1620)) <= "01110110011100000111100001100001";
    rom_arr(integer(1619)) <= "01110010100100100111000011000011";
    rom_arr(integer(1618)) <= "01111010011111101001100001110110";
    rom_arr(integer(1617)) <= "10010011100100111001011110000100";
    rom_arr(integer(1616)) <= "01110100011001110110101001110001";
    rom_arr(integer(1615)) <= "01101110011101100110111110001111";
    rom_arr(integer(1614)) <= "10011000011100100111000001110010";
    rom_arr(integer(1613)) <= "01110000011100110111001001100100";
    rom_arr(integer(1612)) <= "10000001100110110111010010001011";
    rom_arr(integer(1611)) <= "10001001100011101000100110010001";
    rom_arr(integer(1610)) <= "01110101011101111000100001100010";
    rom_arr(integer(1609)) <= "01100111011001100110011001101101";
    rom_arr(integer(1608)) <= "01110010100000010111000010001010";
    rom_arr(integer(1607)) <= "10010100011101010111000001110111";
    rom_arr(integer(1606)) <= "01110010011100100111000101011000";
    rom_arr(integer(1605)) <= "01101100101011111000000010101001";
    rom_arr(integer(1604)) <= "10001111011111111000100010010110";
    rom_arr(integer(1603)) <= "10100010100110010110100101101010";
    rom_arr(integer(1602)) <= "01100100011100111000001010001100";
    rom_arr(integer(1601)) <= "10011000100100011000101110101001";
    rom_arr(integer(1600)) <= "10000101011101010111011101110010";
    rom_arr(integer(1599)) <= "01110001011100010110111101011110";
    rom_arr(integer(1598)) <= "01100010101010001000001101111110";
    rom_arr(integer(1597)) <= "10000100100111110111111010001000";
    rom_arr(integer(1596)) <= "01111010100000101000000110000101";
    rom_arr(integer(1595)) <= "01111001100011110110110101110001";
    rom_arr(integer(1594)) <= "01111001011101010111111110010101";
    rom_arr(integer(1593)) <= "01111011011100110111010001110110";
    rom_arr(integer(1592)) <= "01110001011101010110111101110000";
    rom_arr(integer(1591)) <= "01110011011011100110100001111111";
    rom_arr(integer(1590)) <= "10001000011010101000101101111000";
    rom_arr(integer(1589)) <= "10000111100101100111000110001010";
    rom_arr(integer(1588)) <= "01110101011101111000011010010010";
    rom_arr(integer(1587)) <= "10001010100010011001101010001010";
    rom_arr(integer(1586)) <= "10000000011101010111101001110011";
    rom_arr(integer(1585)) <= "01110010011101110111010101110011";
    rom_arr(integer(1584)) <= "01111001011110111000110110000101";
    rom_arr(integer(1583)) <= "01101000101001010111000110001100";
    rom_arr(integer(1582)) <= "10000101011101101010000101110111";
    rom_arr(integer(1581)) <= "10000111100101111001011110000010";
    rom_arr(integer(1580)) <= "01111001100010011000001010000001";
    rom_arr(integer(1579)) <= "10000100011101010111010001110001";
    rom_arr(integer(1578)) <= "01110010011110000111010001101110";
    rom_arr(integer(1577)) <= "01101111011101100111010101110110";
    rom_arr(integer(1576)) <= "10011111011111000111001110100011";
    rom_arr(integer(1575)) <= "10000110011111001000100010010000";
    rom_arr(integer(1574)) <= "10010001100010101000011101111111";
    rom_arr(integer(1573)) <= "10001110100101011001101010010000";
    rom_arr(integer(1572)) <= "01111101011110010111100101110101";
    rom_arr(integer(1571)) <= "01110001011101100111001001101111";
    rom_arr(integer(1570)) <= "01100100011101000111010101110110";
    rom_arr(integer(1569)) <= "10010001101010101000100010111111";
    rom_arr(integer(1568)) <= "10011111100110101010100010101100";
    rom_arr(integer(1567)) <= "10101001101001011000111110010100";
    rom_arr(integer(1566)) <= "10001011100010111000110101111001";
    rom_arr(integer(1565)) <= "01110111011100010111010101111000";
    rom_arr(integer(1564)) <= "01110100011101000111011101110111";
    rom_arr(integer(1563)) <= "01110000011010100111000110011101";
    rom_arr(integer(1562)) <= "10010010100100111001100110011001";
    rom_arr(integer(1561)) <= "10011000101100111000110010101000";
    rom_arr(integer(1560)) <= "10011110100100001000000110001100";
    rom_arr(integer(1559)) <= "10000001100000101000010001110111";
    rom_arr(integer(1558)) <= "01110001011110010111001001110010";
    rom_arr(integer(1557)) <= "01110111011100100111010101110010";
    rom_arr(integer(1556)) <= "01110101011101010111000101111000";
    rom_arr(integer(1555)) <= "01110001011011110111000001110000";
    rom_arr(integer(1554)) <= "01101101011100100111010101111101";
    rom_arr(integer(1553)) <= "01110111011100010111010101110100";
    rom_arr(integer(1552)) <= "01110100011101100111100001110001";
    rom_arr(integer(1551)) <= "01110001011100110111100001111000";
    rom_arr(integer(1550)) <= "01110111011110000111100101110011";
    rom_arr(integer(1549)) <= "01110111011101010111001001110001";
    rom_arr(integer(1548)) <= "01110011011101110111000101110100";
    rom_arr(integer(1547)) <= "01111001011100100111001101110010";
    rom_arr(integer(1546)) <= "01110010011110010111001001110011";
    rom_arr(integer(1545)) <= "01110110011110010111001001110011";
    rom_arr(integer(1544)) <= "01110110011110100111100001111001";
    rom_arr(integer(1543)) <= "01111000011100110111011001111001";
    rom_arr(integer(1542)) <= "01110110011100110111100001110011";
    rom_arr(integer(1541)) <= "01110111011101010111001001110100";
    rom_arr(integer(1540)) <= "01111001011100110111100101110111";
    rom_arr(integer(1539)) <= "01111001011101100111011001110001";
    rom_arr(integer(1538)) <= "01110110011100100111001001110000";
    rom_arr(integer(1537)) <= "01110101011101000111000101110100";
    rom_arr(integer(1536)) <= "01010011000000000000000000000000";
    rom_arr(integer(1476)) <= "01110101011100010111001001110111";
    rom_arr(integer(1475)) <= "01110101011100000110110101110101";
    rom_arr(integer(1474)) <= "01110101011011110111001001110011";
    rom_arr(integer(1473)) <= "01101111011001100111011001101110";
    rom_arr(integer(1472)) <= "01110010011100010111011001101111";
    rom_arr(integer(1471)) <= "01110010011011110111100001111000";
    rom_arr(integer(1470)) <= "01110100011101000111011101110100";
    rom_arr(integer(1469)) <= "01111000011110000111000101110110";
    rom_arr(integer(1468)) <= "01110101011010100110011001100110";
    rom_arr(integer(1467)) <= "01011010010101000101100101011001";
    rom_arr(integer(1466)) <= "01010111010011100101100101100011";
    rom_arr(integer(1465)) <= "01011110010111100101110101100100";
    rom_arr(integer(1464)) <= "01100111011100000111010101111010";
    rom_arr(integer(1463)) <= "01110001011101000111010001110011";
    rom_arr(integer(1462)) <= "01110011011101000111000001110001";
    rom_arr(integer(1461)) <= "01110001011100000110010101101010";
    rom_arr(integer(1460)) <= "01100010011100100111001001110011";
    rom_arr(integer(1459)) <= "10000110100000101000001001110001";
    rom_arr(integer(1458)) <= "01110111100001100111000101100101";
    rom_arr(integer(1457)) <= "01100111011010110111001101111000";
    rom_arr(integer(1456)) <= "01110111011101000111100101110111";
    rom_arr(integer(1455)) <= "01110110011101010111100101110011";
    rom_arr(integer(1454)) <= "01110011011110000111101101111000";
    rom_arr(integer(1453)) <= "10000011011110010111010010001000";
    rom_arr(integer(1452)) <= "01110010100000110111011101110000";
    rom_arr(integer(1451)) <= "10110111011100111000101101111000";
    rom_arr(integer(1450)) <= "01111011011110010111001101110000";
    rom_arr(integer(1449)) <= "01110100011110000111011001110010";
    rom_arr(integer(1448)) <= "01111000011110010111010101101111";
    rom_arr(integer(1447)) <= "01100111011010101000100110001000";
    rom_arr(integer(1446)) <= "10001011100100110111101010001100";
    rom_arr(integer(1445)) <= "01110001011110110111000101101110";
    rom_arr(integer(1444)) <= "01110001011101101000001110000011";
    rom_arr(integer(1443)) <= "01111100011111000110101001110100";
    rom_arr(integer(1442)) <= "01110001011110010111011101110010";
    rom_arr(integer(1441)) <= "01110010011110000110111101101111";
    rom_arr(integer(1440)) <= "01110001100000111001010001111001";
    rom_arr(integer(1439)) <= "10011101011101110111111001101110";
    rom_arr(integer(1438)) <= "01101011011011000111000001101000";
    rom_arr(integer(1437)) <= "01101111011011110110110101110010";
    rom_arr(integer(1436)) <= "01101101011010100110011101101101";
    rom_arr(integer(1435)) <= "01110010011110100111100101111000";
    rom_arr(integer(1434)) <= "01110111011110000110101101101101";
    rom_arr(integer(1433)) <= "01110111011110110111111010000111";
    rom_arr(integer(1432)) <= "10000010011101101000010001100111";
    rom_arr(integer(1431)) <= "01111011011011010110011101110000";
    rom_arr(integer(1430)) <= "01110110011100110111100110001101";
    rom_arr(integer(1429)) <= "01101000011001000111010001101110";
    rom_arr(integer(1428)) <= "01101111011101110111000101110001";
    rom_arr(integer(1427)) <= "01111000011101100110100101100101";
    rom_arr(integer(1426)) <= "01100001011010110111101001110011";
    rom_arr(integer(1425)) <= "01110001011111101000101110001111";
    rom_arr(integer(1424)) <= "01110111011100010110010001101111";
    rom_arr(integer(1423)) <= "01110101011010100111000101101001";
    rom_arr(integer(1422)) <= "01101010011100100110100001111001";
    rom_arr(integer(1421)) <= "01111100011110000111010101110110";
    rom_arr(integer(1420)) <= "01110010011100110110100001100101";
    rom_arr(integer(1419)) <= "01011101010110011000000001101111";
    rom_arr(integer(1418)) <= "01110001011101010110111001110110";
    rom_arr(integer(1417)) <= "01110101100100000110101101011110";
    rom_arr(integer(1416)) <= "01110111011010110110101001101100";
    rom_arr(integer(1415)) <= "01111000100011101000100101110101";
    rom_arr(integer(1414)) <= "01111110011100000111011001110010";
    rom_arr(integer(1413)) <= "01110010011101010101110101100010";
    rom_arr(integer(1412)) <= "01101110011000101000011110000011";
    rom_arr(integer(1411)) <= "01110111011100010110101010010010";
    rom_arr(integer(1410)) <= "10000000100001101001100010100010";
    rom_arr(integer(1409)) <= "01110101011011001000110110001010";
    rom_arr(integer(1408)) <= "10001000100001000111110101111010";
    rom_arr(integer(1407)) <= "01101100011110000111001001110110";
    rom_arr(integer(1406)) <= "01101111011011100101111101100001";
    rom_arr(integer(1405)) <= "01110011011101001001000101111100";
    rom_arr(integer(1404)) <= "01101011100110001000111110001111";
    rom_arr(integer(1403)) <= "10001100101001000111111101110111";
    rom_arr(integer(1402)) <= "01111110100001111000111010010010";
    rom_arr(integer(1401)) <= "10001111011110100111010001101011";
    rom_arr(integer(1400)) <= "01011100011101000111100101111001";
    rom_arr(integer(1399)) <= "01110100011010000110100101100101";
    rom_arr(integer(1398)) <= "01111010011110011000111110011100";
    rom_arr(integer(1397)) <= "10000011100000111001001110001111";
    rom_arr(integer(1396)) <= "10100011100011110111111010001010";
    rom_arr(integer(1395)) <= "01111100011111111000011110010111";
    rom_arr(integer(1394)) <= "10010111100000100111000101011010";
    rom_arr(integer(1393)) <= "01101001011100010111011101110110";
    rom_arr(integer(1392)) <= "01110000011100110110010101001000";
    rom_arr(integer(1391)) <= "01111011100110100111010101110000";
    rom_arr(integer(1390)) <= "10010001011111111010000110100001";
    rom_arr(integer(1389)) <= "10001001100001000110011110001000";
    rom_arr(integer(1388)) <= "10100001100011111001100010010000";
    rom_arr(integer(1387)) <= "10010011100100101000010010001111";
    rom_arr(integer(1386)) <= "01111110011110100111100101110100";
    rom_arr(integer(1385)) <= "01111000011010000111001001101000";
    rom_arr(integer(1384)) <= "01110011100011001000010010000110";
    rom_arr(integer(1383)) <= "10100101100000001010001010010100";
    rom_arr(integer(1382)) <= "10000111100000010110101110101111";
    rom_arr(integer(1381)) <= "10010011100010011000011110000110";
    rom_arr(integer(1380)) <= "10011000100100111010001010011111";
    rom_arr(integer(1379)) <= "01101111011011000111011001111000";
    rom_arr(integer(1378)) <= "01101111011101000111000101100100";
    rom_arr(integer(1377)) <= "01110100100101001010010010011011";
    rom_arr(integer(1376)) <= "01111111100011001000101010001101";
    rom_arr(integer(1375)) <= "10100100011101100110110010101101";
    rom_arr(integer(1374)) <= "10100100101000011001110010001100";
    rom_arr(integer(1373)) <= "10011010100111101000100101110101";
    rom_arr(integer(1372)) <= "01101000011011100111010101110110";
    rom_arr(integer(1371)) <= "01110100011010110110110001110110";
    rom_arr(integer(1370)) <= "01101111100011101010100110001100";
    rom_arr(integer(1369)) <= "10001000011110110111100010001111";
    rom_arr(integer(1368)) <= "10000110011001110111011011011101";
    rom_arr(integer(1367)) <= "10011101101001110111110010101011";
    rom_arr(integer(1366)) <= "10110000100100101000000101011111";
    rom_arr(integer(1365)) <= "01100011011001100111001101111000";
    rom_arr(integer(1364)) <= "01110101011100100110001101010101";
    rom_arr(integer(1363)) <= "01011100011101000110111001110110";
    rom_arr(integer(1362)) <= "01111101100000001000111110100011";
    rom_arr(integer(1361)) <= "10100101010101100100110010110110";
    rom_arr(integer(1360)) <= "01111011101101001010101110010001";
    rom_arr(integer(1359)) <= "10001110100011111000000001100100";
    rom_arr(integer(1358)) <= "01101111011011000110111101111001";
    rom_arr(integer(1357)) <= "01110100011011110110011001101010";
    rom_arr(integer(1356)) <= "01100011100001101000101101110111";
    rom_arr(integer(1355)) <= "10010001011111110111111101100110";
    rom_arr(integer(1354)) <= "01101111010100010110010110010001";
    rom_arr(integer(1353)) <= "01111100011100111000100101111001";
    rom_arr(integer(1352)) <= "01111001011011010110011101101000";
    rom_arr(integer(1351)) <= "01101001011011110111001001111000";
    rom_arr(integer(1350)) <= "01110001011100100111000001101101";
    rom_arr(integer(1349)) <= "10000111011111101000100010000111";
    rom_arr(integer(1348)) <= "01111011100011010111100110001001";
    rom_arr(integer(1347)) <= "01101010010111010110111101101110";
    rom_arr(integer(1346)) <= "01111011011011100111010101111111";
    rom_arr(integer(1345)) <= "01111010011110000111111001101000";
    rom_arr(integer(1344)) <= "01101100011101100111011001110010";
    rom_arr(integer(1343)) <= "01110110011100001000111010001101";
    rom_arr(integer(1342)) <= "10001011011010001000100101110110";
    rom_arr(integer(1341)) <= "01110000100000000111001001100111";
    rom_arr(integer(1340)) <= "01101010011001010110100001101011";
    rom_arr(integer(1339)) <= "01111111011011111000100001110001";
    rom_arr(integer(1338)) <= "10001010100001111001000001111001";
    rom_arr(integer(1337)) <= "01110101011111000111010101110010";
    rom_arr(integer(1336)) <= "01110110011110110111101110001100";
    rom_arr(integer(1335)) <= "10011011100011101000010001111111";
    rom_arr(integer(1334)) <= "01111101011100110111011101100101";
    rom_arr(integer(1333)) <= "01100111011000100110100001100011";
    rom_arr(integer(1332)) <= "01110100011011101000001101111110";
    rom_arr(integer(1331)) <= "10000110100001001001000110000010";
    rom_arr(integer(1330)) <= "01110011011100100111000001110010";
    rom_arr(integer(1329)) <= "01111001011110100111000101111101";
    rom_arr(integer(1328)) <= "10011101100000000111001101110100";
    rom_arr(integer(1327)) <= "01110100011010000110111001100111";
    rom_arr(integer(1326)) <= "01100000011001110110100001101111";
    rom_arr(integer(1325)) <= "01110010011100101000100001111101";
    rom_arr(integer(1324)) <= "01111100011111001000110001111101";
    rom_arr(integer(1323)) <= "01101110011100100111100001111000";
    rom_arr(integer(1322)) <= "01110100011011100111001101111101";
    rom_arr(integer(1321)) <= "10011001100010100111110110000011";
    rom_arr(integer(1320)) <= "10001011100010010111111110001011";
    rom_arr(integer(1319)) <= "01111101011111010110100110010000";
    rom_arr(integer(1318)) <= "10000111011110111000001001111000";
    rom_arr(integer(1317)) <= "01110100011100000111110001111110";
    rom_arr(integer(1316)) <= "01111001011110000111001001110011";
    rom_arr(integer(1315)) <= "01111001011100100111011010001110";
    rom_arr(integer(1314)) <= "10010010100111111001111110011101";
    rom_arr(integer(1313)) <= "10010011011101111000000010000010";
    rom_arr(integer(1312)) <= "01110100011101010111110101110100";
    rom_arr(integer(1311)) <= "01101111011000110110011001100010";
    rom_arr(integer(1310)) <= "01110001011001100111011101111000";
    rom_arr(integer(1309)) <= "01111001011100100111010101110111";
    rom_arr(integer(1308)) <= "01110001011101100111100101110001";
    rom_arr(integer(1307)) <= "01110110011101010111001101110111";
    rom_arr(integer(1306)) <= "01110010011001100110100101100001";
    rom_arr(integer(1305)) <= "01100000010110010011111001001110";
    rom_arr(integer(1304)) <= "01011000010110100101010001010111";
    rom_arr(integer(1303)) <= "01101011011011110111011101110011";
    rom_arr(integer(1302)) <= "01110100011100110111001101110011";
    rom_arr(integer(1301)) <= "01110001011100010111100101111000";
    rom_arr(integer(1300)) <= "01101111011011100110111001101100";
    rom_arr(integer(1299)) <= "01101111011010100110111001100100";
    rom_arr(integer(1298)) <= "01100101011010100110001101011000";
    rom_arr(integer(1297)) <= "01011110010111100110101101100110";
    rom_arr(integer(1296)) <= "01100110011100000111100001110110";
    rom_arr(integer(1295)) <= "01110110011110010111010001110010";
    rom_arr(integer(1294)) <= "01111001011100100111011101111001";
    rom_arr(integer(1293)) <= "01110101011100000111000101110011";
    rom_arr(integer(1292)) <= "01110101011100100110111101101000";
    rom_arr(integer(1291)) <= "01100011011101010110110101100011";
    rom_arr(integer(1290)) <= "01101001011100100111001101101100";
    rom_arr(integer(1289)) <= "01100111011011100111010101110110";
    rom_arr(integer(1288)) <= "01110001011101100111100101110100";
    rom_arr(integer(1287)) <= "01110001011101010111011101111010";
    rom_arr(integer(1286)) <= "01110100011101000111100001111001";
    rom_arr(integer(1285)) <= "01111000011100010111010101110001";
    rom_arr(integer(1284)) <= "01111000011101010111000101111000";
    rom_arr(integer(1283)) <= "01110111011110010111001101110011";
    rom_arr(integer(1282)) <= "01110110011110010111100101111000";
    rom_arr(integer(1281)) <= "01111001011101000111001001110011";
    rom_arr(integer(1280)) <= "10001001000000000000000000000000";
    rom_arr(integer(1220)) <= "01110010011100010111010101110010";
    rom_arr(integer(1219)) <= "01110011011101100111011101110100";
    rom_arr(integer(1218)) <= "01110100011101010111011101110010";
    rom_arr(integer(1217)) <= "01110010011100110111000101111001";
    rom_arr(integer(1216)) <= "01110010011101100111000101110010";
    rom_arr(integer(1215)) <= "01110110011101000111010001110001";
    rom_arr(integer(1214)) <= "01110110011110010111001101110111";
    rom_arr(integer(1213)) <= "01110101011101010111001001110111";
    rom_arr(integer(1212)) <= "01110111011100110111011101111010";
    rom_arr(integer(1211)) <= "01110010011010010111000001111011";
    rom_arr(integer(1210)) <= "10001011011111010111111110001100";
    rom_arr(integer(1209)) <= "10000001011101010110100001100101";
    rom_arr(integer(1208)) <= "01100111011011010111011001110110";
    rom_arr(integer(1207)) <= "01110111011110010111011101110101";
    rom_arr(integer(1206)) <= "01110001011101000111011110000001";
    rom_arr(integer(1205)) <= "10001011100011011000111010000001";
    rom_arr(integer(1204)) <= "10001100100101011010000110101111";
    rom_arr(integer(1203)) <= "10111000011111111011000110101010";
    rom_arr(integer(1202)) <= "10101011100111101001111001111000";
    rom_arr(integer(1201)) <= "01111001011111010111010110000001";
    rom_arr(integer(1200)) <= "01111001011110010111011001110101";
    rom_arr(integer(1199)) <= "01110100011110100111000101111010";
    rom_arr(integer(1198)) <= "01111111100010110111011010001001";
    rom_arr(integer(1197)) <= "10000001101000101010110110000000";
    rom_arr(integer(1196)) <= "10100001101000011010011110001101";
    rom_arr(integer(1195)) <= "10001011100001111010011110001010";
    rom_arr(integer(1194)) <= "01111011011111000111110101111011";
    rom_arr(integer(1193)) <= "01111001011101010111011001110100";
    rom_arr(integer(1192)) <= "01110011011101000111100010000000";
    rom_arr(integer(1191)) <= "10000101100000000111100110001101";
    rom_arr(integer(1190)) <= "01110111011011110111011110001011";
    rom_arr(integer(1189)) <= "01110010100000110111001010000110";
    rom_arr(integer(1188)) <= "10000001101001000111011110011001";
    rom_arr(integer(1187)) <= "01101101100001111001000010000111";
    rom_arr(integer(1186)) <= "01111111011110000111011101111000";
    rom_arr(integer(1185)) <= "01110110011101001000000010001011";
    rom_arr(integer(1184)) <= "10010010100010110111101110000101";
    rom_arr(integer(1183)) <= "10001101100110100111011110000111";
    rom_arr(integer(1182)) <= "01111110100010001000000010000000";
    rom_arr(integer(1181)) <= "01111110011100010111111101111011";
    rom_arr(integer(1180)) <= "10000011011100010110110110010100";
    rom_arr(integer(1179)) <= "01111010011100100111100001111001";
    rom_arr(integer(1178)) <= "01110100011101000111110010000100";
    rom_arr(integer(1177)) <= "10000111100110111001101010011110";
    rom_arr(integer(1176)) <= "01111110100000001000110001110010";
    rom_arr(integer(1175)) <= "01111110100000100111101001111100";
    rom_arr(integer(1174)) <= "10001011011111101000010010001001";
    rom_arr(integer(1173)) <= "10100100100100100111101110010000";
    rom_arr(integer(1172)) <= "01111001011100000111001101110100";
    rom_arr(integer(1171)) <= "01111001011100111000000001111100";
    rom_arr(integer(1170)) <= "10000111101011000111110001111111";
    rom_arr(integer(1169)) <= "10010110100010011000111110001011";
    rom_arr(integer(1168)) <= "01110101011100111000100001111000";
    rom_arr(integer(1167)) <= "10001010100000001010000110010110";
    rom_arr(integer(1166)) <= "01111000100100011010011101111111";
    rom_arr(integer(1165)) <= "10000010100000000111010101111000";
    rom_arr(integer(1164)) <= "01110100011100010111000110001001";
    rom_arr(integer(1163)) <= "10010101100000101001001010011100";
    rom_arr(integer(1162)) <= "01110011100010000111001001110000";
    rom_arr(integer(1161)) <= "01111101011011101000100110000000";
    rom_arr(integer(1160)) <= "10000110100011100111010010101000";
    rom_arr(integer(1159)) <= "01110110100110100111010010100101";
    rom_arr(integer(1158)) <= "01111100011111100111010101110110";
    rom_arr(integer(1157)) <= "01110110011011110110100110001110";
    rom_arr(integer(1156)) <= "10010000100011000111011101110001";
    rom_arr(integer(1155)) <= "10000001011010011000100101111111";
    rom_arr(integer(1154)) <= "01111111011111110111100101110011";
    rom_arr(integer(1153)) <= "01111110011110110111010101110101";
    rom_arr(integer(1152)) <= "10010010101101101001000110100111";
    rom_arr(integer(1151)) <= "01111011011101110111100001111001";
    rom_arr(integer(1150)) <= "01110101011100000110010001111010";
    rom_arr(integer(1149)) <= "10001100011100001000010001111111";
    rom_arr(integer(1148)) <= "01111111100110101001000101111111";
    rom_arr(integer(1147)) <= "01111000011010010110100001100111";
    rom_arr(integer(1146)) <= "01110001011101010111011101110100";
    rom_arr(integer(1145)) <= "01101101101001111000100101111101";
    rom_arr(integer(1144)) <= "01111010011010110111001001111001";
    rom_arr(integer(1143)) <= "01110000011010110110101101111101";
    rom_arr(integer(1142)) <= "10001111101001010111100110011001";
    rom_arr(integer(1141)) <= "10000000011001100111100101101000";
    rom_arr(integer(1140)) <= "01111010011011110111101101111011";
    rom_arr(integer(1139)) <= "01110110100000000110100001110000";
    rom_arr(integer(1138)) <= "01101000011011110111001001101111";
    rom_arr(integer(1137)) <= "01110100011100110111011101110101";
    rom_arr(integer(1136)) <= "01101110011011010110011010010010";
    rom_arr(integer(1135)) <= "10001101011001011000100101110111";
    rom_arr(integer(1134)) <= "01111001100111010111000101111010";
    rom_arr(integer(1133)) <= "01101101011011100111110010001110";
    rom_arr(integer(1132)) <= "10000010100001111000111001111001";
    rom_arr(integer(1131)) <= "01101111011110110110111101110011";
    rom_arr(integer(1130)) <= "01101111011100110111100101111000";
    rom_arr(integer(1129)) <= "01110100011100100101100101110111";
    rom_arr(integer(1128)) <= "01110100100010100111000101111100";
    rom_arr(integer(1127)) <= "01100111011010010110100101110000";
    rom_arr(integer(1126)) <= "01110111011111010111111010001010";
    rom_arr(integer(1125)) <= "10000001100110011000000010000000";
    rom_arr(integer(1124)) <= "10000001011101010111001110000000";
    rom_arr(integer(1123)) <= "01110101011101010111001001110111";
    rom_arr(integer(1122)) <= "01110011011100110101111100111000";
    rom_arr(integer(1121)) <= "01011001011011010110111110000111";
    rom_arr(integer(1120)) <= "10000011011100110111001001100101";
    rom_arr(integer(1119)) <= "01101011011101111001101010101000";
    rom_arr(integer(1118)) <= "10010110100000010111111101111010";
    rom_arr(integer(1117)) <= "10100001011100101001011110000100";
    rom_arr(integer(1116)) <= "01110010011101000111010101110001";
    rom_arr(integer(1115)) <= "01110101100011000111010100101011";
    rom_arr(integer(1114)) <= "00111110010101000101111101101111";
    rom_arr(integer(1113)) <= "01100111011010010110010001101100";
    rom_arr(integer(1112)) <= "10001000011101001001011110001111";
    rom_arr(integer(1111)) <= "10001110101000010111110110000100";
    rom_arr(integer(1110)) <= "10001110101001010111010101110111";
    rom_arr(integer(1109)) <= "01101100011101110111011101110100";
    rom_arr(integer(1108)) <= "01110001100010111101001011000101";
    rom_arr(integer(1107)) <= "01110011010111000110100001100111";
    rom_arr(integer(1106)) <= "01101001011100100110111101110100";
    rom_arr(integer(1105)) <= "01110010100001101010111010001011";
    rom_arr(integer(1104)) <= "10001011100001001000100110010010";
    rom_arr(integer(1103)) <= "10010000100101100111011001110100";
    rom_arr(integer(1102)) <= "01100010011101000111100101111010";
    rom_arr(integer(1101)) <= "01111010100101011110000011110011";
    rom_arr(integer(1100)) <= "10111110011010010111001001110000";
    rom_arr(integer(1099)) <= "01101111011010100110100001101101";
    rom_arr(integer(1098)) <= "01110100011110101000011010011000";
    rom_arr(integer(1097)) <= "10000110100101011010000110011100";
    rom_arr(integer(1096)) <= "10010100011011100111001001110000";
    rom_arr(integer(1095)) <= "01100111011101000111011101111000";
    rom_arr(integer(1094)) <= "01110111100010111011101111010111";
    rom_arr(integer(1093)) <= "10011000100111111011011001110101";
    rom_arr(integer(1092)) <= "01110101100000110111100101100111";
    rom_arr(integer(1091)) <= "01100110011100000111001001111111";
    rom_arr(integer(1090)) <= "10010001011111100110110001111100";
    rom_arr(integer(1089)) <= "01110100100000010110111001010100";
    rom_arr(integer(1088)) <= "01100010011100000111001001110011";
    rom_arr(integer(1087)) <= "01110101100010001011001111000110";
    rom_arr(integer(1086)) <= "10110001011100111000100010010111";
    rom_arr(integer(1085)) <= "10001100011110011000000001111110";
    rom_arr(integer(1084)) <= "01110000011100110111001101111000";
    rom_arr(integer(1083)) <= "10000000100000111000100101111110";
    rom_arr(integer(1082)) <= "01101101011110100110101001000010";
    rom_arr(integer(1081)) <= "01100101011110000111000101110111";
    rom_arr(integer(1080)) <= "01111000011111101010110010101011";
    rom_arr(integer(1079)) <= "10010111100101011000100001111110";
    rom_arr(integer(1078)) <= "01110101100000110111110110000011";
    rom_arr(integer(1077)) <= "01100100100001110110101010000010";
    rom_arr(integer(1076)) <= "01111101100101100111010010110001";
    rom_arr(integer(1075)) <= "01111001011111000110110001001110";
    rom_arr(integer(1074)) <= "01101000011101010111100101110110";
    rom_arr(integer(1073)) <= "01110110100001001001011110100101";
    rom_arr(integer(1072)) <= "10001011100011110111000110001001";
    rom_arr(integer(1071)) <= "10011010100000010111110101110111";
    rom_arr(integer(1070)) <= "01111000100010110111100010000101";
    rom_arr(integer(1069)) <= "01111000011101100111011001111001";
    rom_arr(integer(1068)) <= "01110111011101010111001001100000";
    rom_arr(integer(1067)) <= "01100110011110010111100101111000";
    rom_arr(integer(1066)) <= "01110010011111011001001010010100";
    rom_arr(integer(1065)) <= "10001100100011100111101010100100";
    rom_arr(integer(1064)) <= "01110100100001011001000110000011";
    rom_arr(integer(1063)) <= "01101100011101011000001001111111";
    rom_arr(integer(1062)) <= "10001000100111110111011001110011";
    rom_arr(integer(1061)) <= "01110100011000100110001001011111";
    rom_arr(integer(1060)) <= "01101111011101000111011001111001";
    rom_arr(integer(1059)) <= "01110011011110001000101110011100";
    rom_arr(integer(1058)) <= "10001110100000011001011101101011";
    rom_arr(integer(1057)) <= "10001011101111101001001010000000";
    rom_arr(integer(1056)) <= "11010111011110000111000110100111";
    rom_arr(integer(1055)) <= "10101001011101010110111101100111";
    rom_arr(integer(1054)) <= "01101110011001010110000101101101";
    rom_arr(integer(1053)) <= "01110010011100100111100001110111";
    rom_arr(integer(1052)) <= "01111001011110100111110001111110";
    rom_arr(integer(1051)) <= "01110001100001011001100010010011";
    rom_arr(integer(1050)) <= "10001000100110001000101001110100";
    rom_arr(integer(1049)) <= "10001111011110100111110101111011";
    rom_arr(integer(1048)) <= "01101101011100000111010001101111";
    rom_arr(integer(1047)) <= "01110010011101100110101101110101";
    rom_arr(integer(1046)) <= "01110110011101110111011101110001";
    rom_arr(integer(1045)) <= "01110011011101010111011001101111";
    rom_arr(integer(1044)) <= "01110010011100010110110001101110";
    rom_arr(integer(1043)) <= "01110111011111100111111001110101";
    rom_arr(integer(1042)) <= "01110000011010110110101001101101";
    rom_arr(integer(1041)) <= "01101011011011000111001101110111";
    rom_arr(integer(1040)) <= "01110110011100110111010101111010";
    rom_arr(integer(1039)) <= "01110100011100110111000101111001";
    rom_arr(integer(1038)) <= "01111010011101100111001001110001";
    rom_arr(integer(1037)) <= "01111000011110000111100001110011";
    rom_arr(integer(1036)) <= "01110001011100100111100001111001";
    rom_arr(integer(1035)) <= "01110110011101100111010001110010";
    rom_arr(integer(1034)) <= "01110010011100010111100001110001";
    rom_arr(integer(1033)) <= "01110001011101100111001001111001";
    rom_arr(integer(1032)) <= "01110100011101110111011101110111";
    rom_arr(integer(1031)) <= "01110111011100100111011101111000";
    rom_arr(integer(1030)) <= "01110011011101000111001001110100";
    rom_arr(integer(1029)) <= "01110101011101110111010001110010";
    rom_arr(integer(1028)) <= "01110100011101000111011101110010";
    rom_arr(integer(1027)) <= "01110010011101000111001101110010";
    rom_arr(integer(1026)) <= "01110101011100010111100101110111";
    rom_arr(integer(1025)) <= "01110101011100010111000001110010";
    rom_arr(integer(1024)) <= "11111110000000000000000000000000";
    rom_arr(integer(964)) <= "01110111011110010111000101110011";
    rom_arr(integer(963)) <= "01110010011100100111010001110100";
    rom_arr(integer(962)) <= "01110011011101100111001101110011";
    rom_arr(integer(961)) <= "01111000011101000111010001111000";
    rom_arr(integer(960)) <= "01110111011101110111000101110101";
    rom_arr(integer(959)) <= "01110100011101110111100001111001";
    rom_arr(integer(958)) <= "01110110011100100111000101110010";
    rom_arr(integer(957)) <= "01110010011110000111000001110001";
    rom_arr(integer(956)) <= "01110001011101000111001001111001";
    rom_arr(integer(955)) <= "01110001011101100111100001111001";
    rom_arr(integer(954)) <= "01110011011101110111001101110010";
    rom_arr(integer(953)) <= "01111000011100010111010001110010";
    rom_arr(integer(952)) <= "01110010011101100111001101110010";
    rom_arr(integer(951)) <= "01111001011110010111010101110011";
    rom_arr(integer(950)) <= "01111000011100010111011001110000";
    rom_arr(integer(949)) <= "01110011011101010111100101110011";
    rom_arr(integer(948)) <= "01101111011100110111001101101111";
    rom_arr(integer(947)) <= "01101010011100000110110101110111";
    rom_arr(integer(946)) <= "01110101011100100111001101110101";
    rom_arr(integer(945)) <= "01110010011101110111000101110110";
    rom_arr(integer(944)) <= "01110110011100100111010101110010";
    rom_arr(integer(943)) <= "01110101011100100111100001110010";
    rom_arr(integer(942)) <= "01110010011100100111000101110000";
    rom_arr(integer(941)) <= "01101101011101010111100101111011";
    rom_arr(integer(940)) <= "01101111011010000110001101100101";
    rom_arr(integer(939)) <= "01011000011000000110010001101010";
    rom_arr(integer(938)) <= "01110010011101000111001101111001";
    rom_arr(integer(937)) <= "01110001011101000111100001110111";
    rom_arr(integer(936)) <= "01110001011110010111001001101101";
    rom_arr(integer(935)) <= "01101101011011100111011010000001";
    rom_arr(integer(934)) <= "10010010100101010111011101110100";
    rom_arr(integer(933)) <= "01110101011110110111010001110110";
    rom_arr(integer(932)) <= "01101111011010010111000001101010";
    rom_arr(integer(931)) <= "01100111011010110111001101110001";
    rom_arr(integer(930)) <= "01111000011101110111011101110000";
    rom_arr(integer(929)) <= "01111001011101100111100001100110";
    rom_arr(integer(928)) <= "01100100011010011000011110001100";
    rom_arr(integer(927)) <= "01111111011110110111011010000101";
    rom_arr(integer(926)) <= "10100111011010011001001010010001";
    rom_arr(integer(925)) <= "01101010100111101000011001111111";
    rom_arr(integer(924)) <= "01110101010111100110011101101011";
    rom_arr(integer(923)) <= "01110101011100110111100001110110";
    rom_arr(integer(922)) <= "01110111011101010110111001110000";
    rom_arr(integer(921)) <= "01101110100000110111001010010111";
    rom_arr(integer(920)) <= "10001111101000111001111110001000";
    rom_arr(integer(919)) <= "10001001100110111001010110100101";
    rom_arr(integer(918)) <= "10001100100011001000101110100111";
    rom_arr(integer(917)) <= "01111100011010100110011001101000";
    rom_arr(integer(916)) <= "01110101011100100111010101110101";
    rom_arr(integer(915)) <= "01110110011101000110110101101101";
    rom_arr(integer(914)) <= "10000000011110001001000110011010";
    rom_arr(integer(913)) <= "01111100100101001000001110001000";
    rom_arr(integer(912)) <= "10001110101000110111111110011111";
    rom_arr(integer(911)) <= "10010100101001101001111101101110";
    rom_arr(integer(910)) <= "10011101011101010111010001101110";
    rom_arr(integer(909)) <= "01110011011101010111100001110111";
    rom_arr(integer(908)) <= "01110011011100100110100001110011";
    rom_arr(integer(907)) <= "10001101100111001000100001111111";
    rom_arr(integer(906)) <= "10000101100001001000101110000011";
    rom_arr(integer(905)) <= "10001011100110011000011110100011";
    rom_arr(integer(904)) <= "10101010101000011001110001111000";
    rom_arr(integer(903)) <= "10001001100100010111100101110011";
    rom_arr(integer(902)) <= "01110010011110100111010101110110";
    rom_arr(integer(901)) <= "01110101011100101000001110000100";
    rom_arr(integer(900)) <= "10001001011101110111110101111010";
    rom_arr(integer(899)) <= "01111001100011001000101110001111";
    rom_arr(integer(898)) <= "01111001011101001001101010110000";
    rom_arr(integer(897)) <= "01111101100011111001000110001001";
    rom_arr(integer(896)) <= "10011110100000000111001001100000";
    rom_arr(integer(895)) <= "01110011011101100111001001110010";
    rom_arr(integer(894)) <= "01110101011010111000101010000110";
    rom_arr(integer(893)) <= "10000111100010111000010110000011";
    rom_arr(integer(892)) <= "10000110100000001000100001110101";
    rom_arr(integer(891)) <= "01110111100100001000100110000101";
    rom_arr(integer(890)) <= "10101100101011011001111110010110";
    rom_arr(integer(889)) <= "10001000100001011000001101011000";
    rom_arr(integer(888)) <= "01110000011101110111100001111000";
    rom_arr(integer(887)) <= "01101111011000111000100010000001";
    rom_arr(integer(886)) <= "01111000100001001000100101111011";
    rom_arr(integer(885)) <= "10001010100010100111001010000001";
    rom_arr(integer(884)) <= "01111101100010000111100001111001";
    rom_arr(integer(883)) <= "10110100100100011001110010001110";
    rom_arr(integer(882)) <= "10010110101001011000010101011011";
    rom_arr(integer(881)) <= "01101000011101010111011101110100";
    rom_arr(integer(880)) <= "01110111011000111000110010000110";
    rom_arr(integer(879)) <= "10000001011110111000110110000110";
    rom_arr(integer(878)) <= "01111010011110101000001001111011";
    rom_arr(integer(877)) <= "01111011100101111000101110010101";
    rom_arr(integer(876)) <= "10010001100010010111111110010001";
    rom_arr(integer(875)) <= "10010000100100000111000001011001";
    rom_arr(integer(874)) <= "01110001011110100111001001111000";
    rom_arr(integer(873)) <= "01110001011001100111111010010000";
    rom_arr(integer(872)) <= "10010001100011111000101001111001";
    rom_arr(integer(871)) <= "01111101011110000110010110001101";
    rom_arr(integer(870)) <= "01111111011100110111100110001011";
    rom_arr(integer(869)) <= "10100100100101101000111110001101";
    rom_arr(integer(868)) <= "01111010100100101000101001011110";
    rom_arr(integer(867)) <= "01110010011100010111011101110101";
    rom_arr(integer(866)) <= "01110010010110100101100110011001";
    rom_arr(integer(865)) <= "10110101100011101001011101111010";
    rom_arr(integer(864)) <= "10000100011100100110110001111101";
    rom_arr(integer(863)) <= "10000100011011111001011010010000";
    rom_arr(integer(862)) <= "01111001100011110111100101110110";
    rom_arr(integer(861)) <= "10001001101010011000100101110001";
    rom_arr(integer(860)) <= "01101111011101010111000101110010";
    rom_arr(integer(859)) <= "01110001010110000110000110011001";
    rom_arr(integer(858)) <= "10111101101001011001001001111001";
    rom_arr(integer(857)) <= "01100011011011010111010001111100";
    rom_arr(integer(856)) <= "01101010011011111001001010010001";
    rom_arr(integer(855)) <= "10100001100001111000111010010011";
    rom_arr(integer(854)) <= "10100010100011010111110001110011";
    rom_arr(integer(853)) <= "01101011011101100111011101110000";
    rom_arr(integer(852)) <= "01110100010110000101001001111000";
    rom_arr(integer(851)) <= "10011011011011101000010101111001";
    rom_arr(integer(850)) <= "01111010011001110110011101110101";
    rom_arr(integer(849)) <= "01011100011101001001011110010001";
    rom_arr(integer(848)) <= "01110111100000101001101110000110";
    rom_arr(integer(847)) <= "10010110011101000111110001110101";
    rom_arr(integer(846)) <= "01110010011100100111100101110100";
    rom_arr(integer(845)) <= "01110011011001100101100001110001";
    rom_arr(integer(844)) <= "01110100011001000111000101110010";
    rom_arr(integer(843)) <= "01101000011001010110011101100100";
    rom_arr(integer(842)) <= "01011100011001110111010001101101";
    rom_arr(integer(841)) <= "01101110011101110110111110000000";
    rom_arr(integer(840)) <= "01111111011100010110110001110010";
    rom_arr(integer(839)) <= "01101011011100110111001101110100";
    rom_arr(integer(838)) <= "01110000011001010101101101101000";
    rom_arr(integer(837)) <= "01101101011011010111101001101110";
    rom_arr(integer(836)) <= "01100100010110100101100101011101";
    rom_arr(integer(835)) <= "01100111011011110101110001101100";
    rom_arr(integer(834)) <= "01110000011001010110101101110000";
    rom_arr(integer(833)) <= "01111100011011100110100110000010";
    rom_arr(integer(832)) <= "01110100011100110111101001111001";
    rom_arr(integer(831)) <= "01101111011011000110010101100001";
    rom_arr(integer(830)) <= "01100101011011010111000101101010";
    rom_arr(integer(829)) <= "01100000010110100110110001101000";
    rom_arr(integer(828)) <= "01011100011000000111010001101001";
    rom_arr(integer(827)) <= "01101111011100000111100001110010";
    rom_arr(integer(826)) <= "01110000011011100111010001110111";
    rom_arr(integer(825)) <= "01101101011101010111010101110101";
    rom_arr(integer(824)) <= "01110101011100110111000010001000";
    rom_arr(integer(823)) <= "01110101011011100111010001101001";
    rom_arr(integer(822)) <= "01101000011010000110101101100111";
    rom_arr(integer(821)) <= "01110001011100110110001101110001";
    rom_arr(integer(820)) <= "01111010011100000111010101110011";
    rom_arr(integer(819)) <= "01111111011000100111011001110011";
    rom_arr(integer(818)) <= "01101111011110000111000101111001";
    rom_arr(integer(817)) <= "01110110011110110111010110001110";
    rom_arr(integer(816)) <= "10001000011100100111010101101111";
    rom_arr(integer(815)) <= "01101000011001100110111101101010";
    rom_arr(integer(814)) <= "01110110011010000110011101110000";
    rom_arr(integer(813)) <= "01101110011010000111010101110111";
    rom_arr(integer(812)) <= "01110101011000110110110001110101";
    rom_arr(integer(811)) <= "01101111011110000111010001111000";
    rom_arr(integer(810)) <= "01111010011101110111001001111111";
    rom_arr(integer(809)) <= "10011110011100101000101010000110";
    rom_arr(integer(808)) <= "10011010100011011000010001110011";
    rom_arr(integer(807)) <= "01101101100000010110110001110101";
    rom_arr(integer(806)) <= "01101011100011110111101110000110";
    rom_arr(integer(805)) <= "01101100011100100110100001110110";
    rom_arr(integer(804)) <= "01101111011100100111010101110110";
    rom_arr(integer(803)) <= "01111010011110000110101101100000";
    rom_arr(integer(802)) <= "10001011100011001000011110000101";
    rom_arr(integer(801)) <= "10000000100000011001000110010011";
    rom_arr(integer(800)) <= "10000010100001011000001101111111";
    rom_arr(integer(799)) <= "01111101100001110111000110000001";
    rom_arr(integer(798)) <= "01110101011111010111100001111011";
    rom_arr(integer(797)) <= "01110100011110010111001001110111";
    rom_arr(integer(796)) <= "01110011011101010110110010000001";
    rom_arr(integer(795)) <= "10001101100001100111111101111001";
    rom_arr(integer(794)) <= "10001101100010000111110110000011";
    rom_arr(integer(793)) <= "10001100100011001001000010001100";
    rom_arr(integer(792)) <= "10010000100011111001000110001000";
    rom_arr(integer(791)) <= "10000111100000010111010001110110";
    rom_arr(integer(790)) <= "01111000011100110111010001110010";
    rom_arr(integer(789)) <= "01110111011110000111000101110110";
    rom_arr(integer(788)) <= "01111110100001101000111110000111";
    rom_arr(integer(787)) <= "10001100100001001000010110000011";
    rom_arr(integer(786)) <= "10000011100010111000101010010011";
    rom_arr(integer(785)) <= "10010100100100111000100110001111";
    rom_arr(integer(784)) <= "10001100011111100111001001111010";
    rom_arr(integer(783)) <= "01110111011100000111000001111001";
    rom_arr(integer(782)) <= "01110111011100100111001001111001";
    rom_arr(integer(781)) <= "01111100011110100111101001111000";
    rom_arr(integer(780)) <= "01111110011111000111011101110101";
    rom_arr(integer(779)) <= "01111000011110001000001010000111";
    rom_arr(integer(778)) <= "01111011011110100111110010000000";
    rom_arr(integer(777)) <= "01111111011111010111100001111001";
    rom_arr(integer(776)) <= "01110001011110010111001101111000";
    rom_arr(integer(775)) <= "01110111011101010111001001110100";
    rom_arr(integer(774)) <= "01111001011110010111000101110110";
    rom_arr(integer(773)) <= "01110100011110010111010101110110";
    rom_arr(integer(772)) <= "01110011011100110111001001111001";
    rom_arr(integer(771)) <= "01110101011100010111000001110110";
    rom_arr(integer(770)) <= "01110010011100100111011001110101";
    rom_arr(integer(769)) <= "01110011011101000111001001110101";
    rom_arr(integer(768)) <= "01101111000000000000000000000000";
    rom_arr(integer(708)) <= "01111001011100110111001101110110";
    rom_arr(integer(707)) <= "01110100100000001000000001111011";
    rom_arr(integer(706)) <= "10000011100001001000000101111111";
    rom_arr(integer(705)) <= "01111100100000011000011001111011";
    rom_arr(integer(704)) <= "01111001011111000111010101111000";
    rom_arr(integer(703)) <= "01110011011101110111000101110010";
    rom_arr(integer(702)) <= "01110111011110100111011001110011";
    rom_arr(integer(701)) <= "01110001011110010111011001110000";
    rom_arr(integer(700)) <= "01110100100000100111100001110110";
    rom_arr(integer(699)) <= "10010110100101101001011110001100";
    rom_arr(integer(698)) <= "10011101100101011001010110000001";
    rom_arr(integer(697)) <= "10000101100011011000110010000100";
    rom_arr(integer(696)) <= "01111011011000100110100001101111";
    rom_arr(integer(695)) <= "01111001011110000111100101110110";
    rom_arr(integer(694)) <= "01110001011110000111011101110001";
    rom_arr(integer(693)) <= "01110001011101010111010101110000";
    rom_arr(integer(692)) <= "01111111100100011001000010011000";
    rom_arr(integer(691)) <= "10011010101000001001100010101110";
    rom_arr(integer(690)) <= "10110110100101111010000110010100";
    rom_arr(integer(689)) <= "10000100011100110111011010000100";
    rom_arr(integer(688)) <= "01110111011101010111010001110111";
    rom_arr(integer(687)) <= "01110100011101100110111101101110";
    rom_arr(integer(686)) <= "01011011011001010110100001101011";
    rom_arr(integer(685)) <= "01101101011010001000010101110011";
    rom_arr(integer(684)) <= "01111001011110111000111101110000";
    rom_arr(integer(683)) <= "01111101100000010111010110001011";
    rom_arr(integer(682)) <= "10001110100101111001101101111111";
    rom_arr(integer(681)) <= "01110111011101010111001101110101";
    rom_arr(integer(680)) <= "01110001011100010111010001101111";
    rom_arr(integer(679)) <= "01010110010101000101000101011001";
    rom_arr(integer(678)) <= "01101000011011010111001001110000";
    rom_arr(integer(677)) <= "01111010011011100110001001100100";
    rom_arr(integer(676)) <= "01100111011011100110111001011101";
    rom_arr(integer(675)) <= "10011100100011110111101001110010";
    rom_arr(integer(674)) <= "01100011011100110111011001111001";
    rom_arr(integer(673)) <= "01110001011100110111010101101111";
    rom_arr(integer(672)) <= "01011001010100010101011101100011";
    rom_arr(integer(671)) <= "01110101011010110110101001110111";
    rom_arr(integer(670)) <= "01110000011101110110000001111101";
    rom_arr(integer(669)) <= "01100111011101010111001001110111";
    rom_arr(integer(668)) <= "10000001011100010111000101011110";
    rom_arr(integer(667)) <= "01100010011010010111010101111010";
    rom_arr(integer(666)) <= "01110110011100110111000001110100";
    rom_arr(integer(665)) <= "01010111010100000101101001100101";
    rom_arr(integer(664)) <= "01100110011010000110100101110100";
    rom_arr(integer(663)) <= "01101000010111110110010001110001";
    rom_arr(integer(662)) <= "01101111011101010110111101110100";
    rom_arr(integer(661)) <= "01011101010111010110001101011010";
    rom_arr(integer(660)) <= "01101000011100000111010101110100";
    rom_arr(integer(659)) <= "01110100011101010110110001101110";
    rom_arr(integer(658)) <= "01100010010100010101111001011010";
    rom_arr(integer(657)) <= "01100111010110100110000101100000";
    rom_arr(integer(656)) <= "01100110011110110111010001111011";
    rom_arr(integer(655)) <= "01101110011011100110111001110011";
    rom_arr(integer(654)) <= "01100110010110110110001001011110";
    rom_arr(integer(653)) <= "01100110011100010111010001110001";
    rom_arr(integer(652)) <= "01110111011110010111010101101111";
    rom_arr(integer(651)) <= "01010101010110100110111001110001";
    rom_arr(integer(650)) <= "01110010011001000110101001101000";
    rom_arr(integer(649)) <= "01101000011111100110111001110100";
    rom_arr(integer(648)) <= "01110001011000000111001101110011";
    rom_arr(integer(647)) <= "01100111011011000110111101110100";
    rom_arr(integer(646)) <= "01101101011111000111011001110110";
    rom_arr(integer(645)) <= "01111001011101010111011101101101";
    rom_arr(integer(644)) <= "01011101011101011000000001110011";
    rom_arr(integer(643)) <= "01110100011101100111011101110010";
    rom_arr(integer(642)) <= "01110001011100101000001101101110";
    rom_arr(integer(641)) <= "01111000011101000110111101101110";
    rom_arr(integer(640)) <= "01101100011001110111111101111101";
    rom_arr(integer(639)) <= "01101110011101110111010001110001";
    rom_arr(integer(638)) <= "01110000011101110111110110000010";
    rom_arr(integer(637)) <= "01110110100000000111010110001100";
    rom_arr(integer(636)) <= "01101110100011010111011001110111";
    rom_arr(integer(635)) <= "10001000100001011000000110000110";
    rom_arr(integer(634)) <= "01101101011001110111001001110100";
    rom_arr(integer(633)) <= "01101111011101011000000010000010";
    rom_arr(integer(632)) <= "01101010011100010111011001110001";
    rom_arr(integer(631)) <= "01110001011011110110011101101000";
    rom_arr(integer(630)) <= "01110010011100101001010110011000";
    rom_arr(integer(629)) <= "10010010011110111001100001111000";
    rom_arr(integer(628)) <= "10001011010110010111110101101110";
    rom_arr(integer(627)) <= "01011010011010000111000001111001";
    rom_arr(integer(626)) <= "10100111011101110110111001111101";
    rom_arr(integer(625)) <= "01101101011101110111001101110100";
    rom_arr(integer(624)) <= "01110010011011100110000001101011";
    rom_arr(integer(623)) <= "10010111101000011000111110010110";
    rom_arr(integer(622)) <= "01111011101000111100000001011111";
    rom_arr(integer(621)) <= "10001100011001100110110001011100";
    rom_arr(integer(620)) <= "01100111011100010110101101101100";
    rom_arr(integer(619)) <= "01110001011110100111001101110000";
    rom_arr(integer(618)) <= "10000011011101110111000001110110";
    rom_arr(integer(617)) <= "01110010011110000110111001110010";
    rom_arr(integer(616)) <= "10010100100010100111000110011111";
    rom_arr(integer(615)) <= "11000011100011011000100110001001";
    rom_arr(integer(614)) <= "01110001011100010110001001011001";
    rom_arr(integer(613)) <= "01100011011101000111000101111010";
    rom_arr(integer(612)) <= "01110110011101101001000110001001";
    rom_arr(integer(611)) <= "10001001100000000111101001110100";
    rom_arr(integer(610)) <= "01110011011101010111110001111010";
    rom_arr(integer(609)) <= "01101100011110011010000010010000";
    rom_arr(integer(608)) <= "01100111011100110111101010001110";
    rom_arr(integer(607)) <= "01111010011100010101100101001111";
    rom_arr(integer(606)) <= "01110000100001100111000001101000";
    rom_arr(integer(605)) <= "10000000101100101000001110001110";
    rom_arr(integer(604)) <= "10011000100010100111011001111000";
    rom_arr(integer(603)) <= "01110011011111010111011001100101";
    rom_arr(integer(602)) <= "01101110101010111000111001111001";
    rom_arr(integer(601)) <= "01111010101000001001011110100111";
    rom_arr(integer(600)) <= "10101011011011010101000001011101";
    rom_arr(integer(599)) <= "10011000011100010111000011011010";
    rom_arr(integer(598)) <= "10101001011110011000100010011110";
    rom_arr(integer(597)) <= "10100000100110010111111001110101";
    rom_arr(integer(596)) <= "01110111011100110110111001100101";
    rom_arr(integer(595)) <= "01110000100111001001001010101010";
    rom_arr(integer(594)) <= "10000010101010011000111110001011";
    rom_arr(integer(593)) <= "10100110101100111000100010000110";
    rom_arr(integer(592)) <= "10010100101101101001000001101110";
    rom_arr(integer(591)) <= "10010001100001100111111010001101";
    rom_arr(integer(590)) <= "10010001100110110111110001110101";
    rom_arr(integer(589)) <= "01110010011110110111011101101011";
    rom_arr(integer(588)) <= "01110111100111001001101010101011";
    rom_arr(integer(587)) <= "10100001100010111000011010110100";
    rom_arr(integer(586)) <= "10001100100010001001100001100111";
    rom_arr(integer(585)) <= "01100110011101101001000101111000";
    rom_arr(integer(584)) <= "10000110100011101000110110001111";
    rom_arr(integer(583)) <= "10010001100010110111111101110010";
    rom_arr(integer(582)) <= "10000000011101010111100001111100";
    rom_arr(integer(581)) <= "10000011100100011001011101110110";
    rom_arr(integer(580)) <= "10010100100101111011010110001111";
    rom_arr(integer(579)) <= "10010100101010010111100110100011";
    rom_arr(integer(578)) <= "10000010011110001000110010000111";
    rom_arr(integer(577)) <= "10000110100100111000101010010001";
    rom_arr(integer(576)) <= "10001111100000000111110101110111";
    rom_arr(integer(575)) <= "01110101011101100110101001110010";
    rom_arr(integer(574)) <= "10001100100100100111010110010101";
    rom_arr(integer(573)) <= "10000010100111101000001010001000";
    rom_arr(integer(572)) <= "10011000100010100110111110011100";
    rom_arr(integer(571)) <= "10010010011111111001000110011000";
    rom_arr(integer(570)) <= "10100101100011101000101110001100";
    rom_arr(integer(569)) <= "10010101100000000111101001110010";
    rom_arr(integer(568)) <= "01110100011110010111001001111000";
    rom_arr(integer(567)) <= "10000000100000111000110110100100";
    rom_arr(integer(566)) <= "01110111101000111000101010001011";
    rom_arr(integer(565)) <= "10001001011011011000110110001111";
    rom_arr(integer(564)) <= "01111011100011101000110101111011";
    rom_arr(integer(563)) <= "10011001100011000111110110001010";
    rom_arr(integer(562)) <= "10010011011111110111010101111001";
    rom_arr(integer(561)) <= "01111000011110000111000101101101";
    rom_arr(integer(560)) <= "01100101011101001000011101110011";
    rom_arr(integer(559)) <= "01111001011111111000101010000101";
    rom_arr(integer(558)) <= "01111100011110110111010010010010";
    rom_arr(integer(557)) <= "10101110100011101000111010011010";
    rom_arr(integer(556)) <= "10010000100101011000110101111111";
    rom_arr(integer(555)) <= "10000110011101000111010001110101";
    rom_arr(integer(554)) <= "01110111011110000111000101110000";
    rom_arr(integer(553)) <= "01101111011010010110011101011011";
    rom_arr(integer(552)) <= "01100101011011100110111001110011";
    rom_arr(integer(551)) <= "01110001011100101000000110001011";
    rom_arr(integer(550)) <= "01110111011101101001010110010010";
    rom_arr(integer(549)) <= "10000100011110100111110001110010";
    rom_arr(integer(548)) <= "01110100011101000111100101110010";
    rom_arr(integer(547)) <= "01110101011101100111011101110001";
    rom_arr(integer(546)) <= "01110100011100010111010101101111";
    rom_arr(integer(545)) <= "01101010011010110110011101100110";
    rom_arr(integer(544)) <= "01100101011001010110100001100100";
    rom_arr(integer(543)) <= "01011100010101110101111101101001";
    rom_arr(integer(542)) <= "01101011011011000111010001110110";
    rom_arr(integer(541)) <= "01110001011100100111001101110101";
    rom_arr(integer(540)) <= "01110111011100110111100101110111";
    rom_arr(integer(539)) <= "01110111011110000111011001110111";
    rom_arr(integer(538)) <= "01110100011101110110111001110001";
    rom_arr(integer(537)) <= "01101101011011110110100101101011";
    rom_arr(integer(536)) <= "01101001011010000111001101110010";
    rom_arr(integer(535)) <= "01110101011101110111101001111000";
    rom_arr(integer(534)) <= "01110100011100010111001101111001";
    rom_arr(integer(533)) <= "01110011011101100111001101110101";
    rom_arr(integer(532)) <= "01110000011110010111001001110001";
    rom_arr(integer(531)) <= "01110010011101100111001001110101";
    rom_arr(integer(530)) <= "01110100011100010111010001110101";
    rom_arr(integer(529)) <= "01110100011100000111000001110111";
    rom_arr(integer(528)) <= "01110101011101110111010001111000";
    rom_arr(integer(527)) <= "01110101011101010111000101111000";
    rom_arr(integer(526)) <= "01110001011110010111100001110001";
    rom_arr(integer(525)) <= "01110001011100110111000101110111";
    rom_arr(integer(524)) <= "01110100011110010111011001110110";
    rom_arr(integer(523)) <= "01110100011110000111000101110100";
    rom_arr(integer(522)) <= "01110111011101110111101001111001";
    rom_arr(integer(521)) <= "01110001011101100111000101111001";
    rom_arr(integer(520)) <= "01111001011101110111100101110011";
    rom_arr(integer(519)) <= "01110011011110010111001001110110";
    rom_arr(integer(518)) <= "01110110011101000111000101110010";
    rom_arr(integer(517)) <= "01110000011101110111001001110001";
    rom_arr(integer(516)) <= "01110111011110000111011101110101";
    rom_arr(integer(515)) <= "01110100011100110111001001110001";
    rom_arr(integer(514)) <= "01110101011110010111000101110100";
    rom_arr(integer(513)) <= "01111001011101000111001101111001";
    rom_arr(integer(512)) <= "11010100000000000000000000000000";
    rom_arr(integer(452)) <= "01111001011110010111100001110111";
    rom_arr(integer(451)) <= "01110011011101100111000101110011";
    rom_arr(integer(450)) <= "01110101011110010111001101110101";
    rom_arr(integer(449)) <= "01110001011101100111100101110101";
    rom_arr(integer(448)) <= "01111001011101010111100001110100";
    rom_arr(integer(447)) <= "01111010011101110111010001110011";
    rom_arr(integer(446)) <= "01110010011110000111101001110011";
    rom_arr(integer(445)) <= "01110110011101100111010001110110";
    rom_arr(integer(444)) <= "01110001011101000111000001101010";
    rom_arr(integer(443)) <= "01101111011100010111000101101010";
    rom_arr(integer(442)) <= "01100111011010110111010001110100";
    rom_arr(integer(441)) <= "01110011011011000111000101110100";
    rom_arr(integer(440)) <= "01110101011010110111010101110111";
    rom_arr(integer(439)) <= "01110110011101110111100001110011";
    rom_arr(integer(438)) <= "01110100011101100111100101110100";
    rom_arr(integer(437)) <= "01101101011100110110111101111011";
    rom_arr(integer(436)) <= "10001001100001011010101110100000";
    rom_arr(integer(435)) <= "10100110101001100111110010001101";
    rom_arr(integer(434)) <= "10101011101001000111000101110000";
    rom_arr(integer(433)) <= "01110001011100000110001001101101";
    rom_arr(integer(432)) <= "01111001011100110111100101110011";
    rom_arr(integer(431)) <= "01110001011100100111010101101100";
    rom_arr(integer(430)) <= "01110001011100000111001010001000";
    rom_arr(integer(429)) <= "10111111100111100110011111001000";
    rom_arr(integer(428)) <= "10001010101010001001001010010101";
    rom_arr(integer(427)) <= "10100011011111011000001110011111";
    rom_arr(integer(426)) <= "01110000011001100101110001100110";
    rom_arr(integer(425)) <= "01101011011101100111011101110110";
    rom_arr(integer(424)) <= "01110101011101010111001001101110";
    rom_arr(integer(423)) <= "10000100100000001000000110001000";
    rom_arr(integer(422)) <= "10010101101000010111101010000110";
    rom_arr(integer(421)) <= "10000101011110111001011110000101";
    rom_arr(integer(420)) <= "10000010011111000111111010011111";
    rom_arr(integer(419)) <= "01101011011010000110101101110100";
    rom_arr(integer(418)) <= "01110100011110010111011001111001";
    rom_arr(integer(417)) <= "01110111011100100111000001101110";
    rom_arr(integer(416)) <= "01111101011110111000101001101011";
    rom_arr(integer(415)) <= "01110100011111110111110001110100";
    rom_arr(integer(414)) <= "01111111100001010111100101111101";
    rom_arr(integer(413)) <= "10000011011110100111100001101110";
    rom_arr(integer(412)) <= "10001010100011010111100001111101";
    rom_arr(integer(411)) <= "01110101011100010111001101110001";
    rom_arr(integer(410)) <= "01110100011101100110111101100010";
    rom_arr(integer(409)) <= "01110110100011110110111110001110";
    rom_arr(integer(408)) <= "01111111011111101001000101110010";
    rom_arr(integer(407)) <= "01110011011101111000001001101000";
    rom_arr(integer(406)) <= "01111101011010111001010101110110";
    rom_arr(integer(405)) <= "10100011101000000111010001110110";
    rom_arr(integer(404)) <= "01101010011101100111011001110101";
    rom_arr(integer(403)) <= "01110111011101100110100101100111";
    rom_arr(integer(402)) <= "10001010100011001011000110011101";
    rom_arr(integer(401)) <= "10001010011110000111100101101010";
    rom_arr(integer(400)) <= "10000010011001011000001001111110";
    rom_arr(integer(399)) <= "01110101100100100111110010001000";
    rom_arr(integer(398)) <= "10101001011110010111011001101111";
    rom_arr(integer(397)) <= "01100110011100010111001101111000";
    rom_arr(integer(396)) <= "01110110011100100110010001101011";
    rom_arr(integer(395)) <= "10100110101000100110101101110100";
    rom_arr(integer(394)) <= "10000000100010001000001101111110";
    rom_arr(integer(393)) <= "01110010011100100111001110000011";
    rom_arr(integer(392)) <= "01110011100011101000111010000011";
    rom_arr(integer(391)) <= "01101111100001101010010001101110";
    rom_arr(integer(390)) <= "01100111011101000111001101110010";
    rom_arr(integer(389)) <= "01111001011101000110001001110001";
    rom_arr(integer(388)) <= "10010000011100110110111110000011";
    rom_arr(integer(387)) <= "01110001011101100110110101110011";
    rom_arr(integer(386)) <= "01110110011101011000010110001101";
    rom_arr(integer(385)) <= "10010111100101101001001101111111";
    rom_arr(integer(384)) <= "01110100100110000111010001101100";
    rom_arr(integer(383)) <= "01101100011101000111010101110011";
    rom_arr(integer(382)) <= "01111000011100000110001010000111";
    rom_arr(integer(381)) <= "10001110011101010111101101110101";
    rom_arr(integer(380)) <= "01110111011001100111011110000110";
    rom_arr(integer(379)) <= "01110000100000111000100110010001";
    rom_arr(integer(378)) <= "10001100100000111001110110001011";
    rom_arr(integer(377)) <= "10110011011100000111000101110010";
    rom_arr(integer(376)) <= "01110101011101100111010101110011";
    rom_arr(integer(375)) <= "01110100011011110110100001101010";
    rom_arr(integer(374)) <= "10000100011011000111000101101101";
    rom_arr(integer(373)) <= "01100111011100111000100010001000";
    rom_arr(integer(372)) <= "01111110100001101000101010011001";
    rom_arr(integer(371)) <= "10000101100100100111110101110101";
    rom_arr(integer(370)) <= "01110100011101010110101101101000";
    rom_arr(integer(369)) <= "01111010011101010111001001110110";
    rom_arr(integer(368)) <= "01110110011100000111101001100101";
    rom_arr(integer(367)) <= "01101010011101000111001101110000";
    rom_arr(integer(366)) <= "01111001100001000111011101111001";
    rom_arr(integer(365)) <= "10000001100110101001000010001101";
    rom_arr(integer(364)) <= "01111001011101011000011001110001";
    rom_arr(integer(363)) <= "01110101011100110110011101101001";
    rom_arr(integer(362)) <= "01110011011101100111010101111001";
    rom_arr(integer(361)) <= "01110011011101010111101101100111";
    rom_arr(integer(360)) <= "01100011011001110111010001101011";
    rom_arr(integer(359)) <= "01111101011101001000001110000010";
    rom_arr(integer(358)) <= "10000011100010101001100110001110";
    rom_arr(integer(357)) <= "10011100100000010110100101101011";
    rom_arr(integer(356)) <= "01101101011110010111100001100101";
    rom_arr(integer(355)) <= "01110111011101000111011101110000";
    rom_arr(integer(354)) <= "01111000011101010111110110010000";
    rom_arr(integer(353)) <= "10011100100010000110101010101100";
    rom_arr(integer(352)) <= "01110110011111010110111110001000";
    rom_arr(integer(351)) <= "10011001011101111010100010011001";
    rom_arr(integer(350)) <= "10010000011011101000000001111110";
    rom_arr(integer(349)) <= "01111011100110001000001001110010";
    rom_arr(integer(348)) <= "01111011011101110111100101110000";
    rom_arr(integer(347)) <= "01110000011101110111100110111100";
    rom_arr(integer(346)) <= "10110001101000011011000110001001";
    rom_arr(integer(345)) <= "10011100011100111000011101111101";
    rom_arr(integer(344)) <= "10000111100001101001111010001101";
    rom_arr(integer(343)) <= "10000111011111001000110001101101";
    rom_arr(integer(342)) <= "10100100011100001010010001111000";
    rom_arr(integer(341)) <= "01111110011110010111011101110100";
    rom_arr(integer(340)) <= "01110101100001100111100110010111";
    rom_arr(integer(339)) <= "10010110100100010111100110000000";
    rom_arr(integer(338)) <= "01110101011010010111000001111001";
    rom_arr(integer(337)) <= "01111110101101001001101010001111";
    rom_arr(integer(336)) <= "10001011100100101010001010100110";
    rom_arr(integer(335)) <= "11000110100010101000111010000001";
    rom_arr(integer(334)) <= "01110001011100010111011001110101";
    rom_arr(integer(333)) <= "01110101011110100111001001110110";
    rom_arr(integer(332)) <= "10010011100100001001001110010000";
    rom_arr(integer(331)) <= "10011101100100110111011001101100";
    rom_arr(integer(330)) <= "01011110011101010111100110011011";
    rom_arr(integer(329)) <= "10000011100110001000100101111010";
    rom_arr(integer(328)) <= "01110101100001000111010010010010";
    rom_arr(integer(327)) <= "01101110011100110111011001110100";
    rom_arr(integer(326)) <= "01110010100100001001011110011100";
    rom_arr(integer(325)) <= "10011010100010011000111010000001";
    rom_arr(integer(324)) <= "10000001011101101000101101111100";
    rom_arr(integer(323)) <= "01100101011101110111110001101001";
    rom_arr(integer(322)) <= "10000111011110001000101110010000";
    rom_arr(integer(321)) <= "01111110100100110111011101110110";
    rom_arr(integer(320)) <= "01110010011101100111010001110110";
    rom_arr(integer(319)) <= "01111111100010011001000110110011";
    rom_arr(integer(318)) <= "10001010100001011000111110000010";
    rom_arr(integer(317)) <= "10010010100010110111011110001111";
    rom_arr(integer(316)) <= "01110011011011101000101110000110";
    rom_arr(integer(315)) <= "01111001100010101000101101110001";
    rom_arr(integer(314)) <= "10011011100101101000100101111001";
    rom_arr(integer(313)) <= "01111100011100110111010001110001";
    rom_arr(integer(312)) <= "01110011011101100111111010011001";
    rom_arr(integer(311)) <= "10101000011111001001010001110010";
    rom_arr(integer(310)) <= "01110111100010000110111001111011";
    rom_arr(integer(309)) <= "10001110011000000111110101101110";
    rom_arr(integer(308)) <= "01101101100001000111001110100111";
    rom_arr(integer(307)) <= "01101100011011100111010101110010";
    rom_arr(integer(306)) <= "01110000011100010111011101110001";
    rom_arr(integer(305)) <= "01110010011101111001001101110001";
    rom_arr(integer(304)) <= "10011101011101010111011110000001";
    rom_arr(integer(303)) <= "10011111011011111000110101111110";
    rom_arr(integer(302)) <= "10001111100000001000000010011011";
    rom_arr(integer(301)) <= "01110101011110101000001001111010";
    rom_arr(integer(300)) <= "01110011011011110110111001101111";
    rom_arr(integer(299)) <= "01110110011100100111011001110100";
    rom_arr(integer(298)) <= "01111000011101101000111010000011";
    rom_arr(integer(297)) <= "01101101011101110111111010010111";
    rom_arr(integer(296)) <= "10001000011011011010000010000111";
    rom_arr(integer(295)) <= "01111111100010011000000010010000";
    rom_arr(integer(294)) <= "10100011011011011000011001110001";
    rom_arr(integer(293)) <= "10000010011011000110101101110101";
    rom_arr(integer(292)) <= "01110000011101100111100001110110";
    rom_arr(integer(291)) <= "01111000011111001000010110000110";
    rom_arr(integer(290)) <= "01111110100100001000000110100111";
    rom_arr(integer(289)) <= "01110010101110011000101110110011";
    rom_arr(integer(288)) <= "10100001110001010110010011011101";
    rom_arr(integer(287)) <= "10001011100111001001000010000101";
    rom_arr(integer(286)) <= "01110010011011000111000101110011";
    rom_arr(integer(285)) <= "01110110011100100111010101110100";
    rom_arr(integer(284)) <= "01111000011100010111010001110101";
    rom_arr(integer(283)) <= "10000010100010000111110101110010";
    rom_arr(integer(282)) <= "01110001100011101000001101110110";
    rom_arr(integer(281)) <= "01110110011101010111100101110011";
    rom_arr(integer(280)) <= "01110100011110010111010101111000";
    rom_arr(integer(279)) <= "01110001011100100111001001110001";
    rom_arr(integer(278)) <= "01110010011101010111100101110110";
    rom_arr(integer(277)) <= "01110011011101000111001001111001";
    rom_arr(integer(276)) <= "01110101011100110111001001110101";
    rom_arr(integer(275)) <= "01110011011101010110111001101110";
    rom_arr(integer(274)) <= "01110000011100110111000101110000";
    rom_arr(integer(273)) <= "01110000011100000111100001110100";
    rom_arr(integer(272)) <= "01110011011110010111000101110110";
    rom_arr(integer(271)) <= "01110110011100100111010101110010";
    rom_arr(integer(270)) <= "01110011011101110111010001111001";
    rom_arr(integer(269)) <= "01110100011100010111011101110011";
    rom_arr(integer(268)) <= "01111000011100010111010101110110";
    rom_arr(integer(267)) <= "01110110011101110111100001110011";
    rom_arr(integer(266)) <= "01110010011101000111100101111000";
    rom_arr(integer(265)) <= "01111010011100100111100101110001";
    rom_arr(integer(264)) <= "01111001011100100111011101111000";
    rom_arr(integer(263)) <= "01110001011100100111001001110011";
    rom_arr(integer(262)) <= "01110010011101000111011001111010";
    rom_arr(integer(261)) <= "01110001011101010111100101111000";
    rom_arr(integer(260)) <= "01110111011101000111011101110101";
    rom_arr(integer(259)) <= "01110110011100000111001001110100";
    rom_arr(integer(258)) <= "01110011011101000111001001111001";
    rom_arr(integer(257)) <= "01111000011101100111000101110001";
    rom_arr(integer(256)) <= "00000000000000000000000000000000";
    rom_arr(integer(196)) <= "01110101011110000111100101110111";
    rom_arr(integer(195)) <= "01111000011101100111100001111000";
    rom_arr(integer(194)) <= "01110000011101000111001001110001";
    rom_arr(integer(193)) <= "01111011011101100110100101111010";
    rom_arr(integer(192)) <= "01110011011101110111011101111000";
    rom_arr(integer(191)) <= "01111001011101100111001101111000";
    rom_arr(integer(190)) <= "01110011011110100111100001110110";
    rom_arr(integer(189)) <= "01111001011101010111010001110111";
    rom_arr(integer(188)) <= "01111010011101111000100010001101";
    rom_arr(integer(187)) <= "10001101101001001001011010011100";
    rom_arr(integer(186)) <= "10010111101110001010010010101111";
    rom_arr(integer(185)) <= "10100001101001011010110010100010";
    rom_arr(integer(184)) <= "10100001100110101000111001111110";
    rom_arr(integer(183)) <= "01110111011100110111001001110110";
    rom_arr(integer(182)) <= "01110011011101000111011001101110";
    rom_arr(integer(181)) <= "01111011011101101001001010011100";
    rom_arr(integer(180)) <= "10001101100100101001010110011101";
    rom_arr(integer(179)) <= "10010011101010101001100110100101";
    rom_arr(integer(178)) <= "10100000101001011001001010011101";
    rom_arr(integer(177)) <= "10010000100100001001110001110111";
    rom_arr(integer(176)) <= "01110001011100010111011001111000";
    rom_arr(integer(175)) <= "01110010011100100111000001101011";
    rom_arr(integer(174)) <= "10001011100011111000011110001111";
    rom_arr(integer(173)) <= "10001001100010001000101010000110";
    rom_arr(integer(172)) <= "10000001011001110111000101110010";
    rom_arr(integer(171)) <= "10000000100010110110101110010001";
    rom_arr(integer(170)) <= "10000011011111000111100101110111";
    rom_arr(integer(169)) <= "01110001011110010111011101110010";
    rom_arr(integer(168)) <= "01110100011100010111010010000101";
    rom_arr(integer(167)) <= "10000110100111001000101001111100";
    rom_arr(integer(166)) <= "01111110011110000111001001110011";
    rom_arr(integer(165)) <= "01101101011111110111000101101111";
    rom_arr(integer(164)) <= "01110000011100100110100010000001";
    rom_arr(integer(163)) <= "01101111011011000110100101100111";
    rom_arr(integer(162)) <= "01110001011101000111000001110010";
    rom_arr(integer(161)) <= "01110110011101100111011110000000";
    rom_arr(integer(160)) <= "10000101011100100110110101111000";
    rom_arr(integer(159)) <= "01101000011011110110111001101100";
    rom_arr(integer(158)) <= "01011101011110010110100001111001";
    rom_arr(integer(157)) <= "01110110100001110110111110001011";
    rom_arr(integer(156)) <= "01110100011100100110011001101110";
    rom_arr(integer(155)) <= "01110110011101100111101001111001";
    rom_arr(integer(154)) <= "01110101011100110111010010000100";
    rom_arr(integer(153)) <= "01110101011010000111011101110100";
    rom_arr(integer(152)) <= "01110100011010110110100001110000";
    rom_arr(integer(151)) <= "01100100010111000101111001100011";
    rom_arr(integer(150)) <= "01100011011011010111000101110001";
    rom_arr(integer(149)) <= "01110100011111100111100001101110";
    rom_arr(integer(148)) <= "01101110011101110111000101110001";
    rom_arr(integer(147)) <= "01111001011101110111101010000100";
    rom_arr(integer(146)) <= "01110100011011110110100001110000";
    rom_arr(integer(145)) <= "01111001011100010111100001110111";
    rom_arr(integer(144)) <= "01100100011011000110101101011001";
    rom_arr(integer(143)) <= "01011011011001110110110001110010";
    rom_arr(integer(142)) <= "01101111011101010111111101101101";
    rom_arr(integer(141)) <= "01100101011100100111000101110001";
    rom_arr(integer(140)) <= "01110011011101000110110101101101";
    rom_arr(integer(139)) <= "01100111011010010111000001111110";
    rom_arr(integer(138)) <= "10000010011101000110011101110101";
    rom_arr(integer(137)) <= "01100100011010000110110001110101";
    rom_arr(integer(136)) <= "01101000011011100110111001111001";
    rom_arr(integer(135)) <= "10001010011111010110100101100011";
    rom_arr(integer(134)) <= "01101000011101000111001001110101";
    rom_arr(integer(133)) <= "01110011011100010110110101010110";
    rom_arr(integer(132)) <= "01011011011011010111010010000011";
    rom_arr(integer(131)) <= "01101111011100100111111101111011";
    rom_arr(integer(130)) <= "01111110100011010110101001101000";
    rom_arr(integer(129)) <= "10010100101010010111000001110001";
    rom_arr(integer(128)) <= "01111101100010010110011101100011";
    rom_arr(integer(127)) <= "01101000011101000111011101110100";
    rom_arr(integer(126)) <= "01110101011101100110110101011001";
    rom_arr(integer(125)) <= "01100001011011110111010001110100";
    rom_arr(integer(124)) <= "01110001011111101000000101111011";
    rom_arr(integer(123)) <= "10010000011101111000010010000111";
    rom_arr(integer(122)) <= "01110000100011000111100110010001";
    rom_arr(integer(121)) <= "10001011011100000111000001100100";
    rom_arr(integer(120)) <= "01101010011100100111100101110101";
    rom_arr(integer(119)) <= "01111010011100110110010001010110";
    rom_arr(integer(118)) <= "01100001100001000111000101111001";
    rom_arr(integer(117)) <= "01101011100000111000111110001011";
    rom_arr(integer(116)) <= "01111010011111000111001101110111";
    rom_arr(integer(115)) <= "10001011100001110111000110001111";
    rom_arr(integer(114)) <= "01111100011101001000001110000001";
    rom_arr(integer(113)) <= "01110000011100000111001101110010";
    rom_arr(integer(112)) <= "01110100011011100110110001010100";
    rom_arr(integer(111)) <= "01100110011110110111000110000100";
    rom_arr(integer(110)) <= "10001100100000001001110110001100";
    rom_arr(integer(109)) <= "10001101011011100111101101110100";
    rom_arr(integer(108)) <= "10001001100000110111101010001000";
    rom_arr(integer(107)) <= "10000010100001000111111010000011";
    rom_arr(integer(106)) <= "01110100011011000111100101111000";
    rom_arr(integer(105)) <= "01110111011100010110100101010001";
    rom_arr(integer(104)) <= "01011110011111101001010010010001";
    rom_arr(integer(103)) <= "01111111100001101001010010001111";
    rom_arr(integer(102)) <= "10001010011111001000111010000001";
    rom_arr(integer(101)) <= "10000000100000110111110101110101";
    rom_arr(integer(100)) <= "10000010101000010111111110010010";
    rom_arr(integer(99)) <= "01110100011100000111011001110100";
    rom_arr(integer(98)) <= "01110110011011000110000001010011";
    rom_arr(integer(97)) <= "01101010100001111001110010011000";
    rom_arr(integer(96)) <= "10011110100010001000101010011110";
    rom_arr(integer(95)) <= "10010001100010011000111101111001";
    rom_arr(integer(94)) <= "10000101100001000111100010001111";
    rom_arr(integer(93)) <= "10100000011111111001001010110011";
    rom_arr(integer(92)) <= "01101110011001110111001001111001";
    rom_arr(integer(91)) <= "01110111011011110110101001100000";
    rom_arr(integer(90)) <= "10100110101001101010101010001000";
    rom_arr(integer(89)) <= "10010101100101011000110010001110";
    rom_arr(integer(88)) <= "10010111100011001000010001110101";
    rom_arr(integer(87)) <= "10010111100100111001011110010111";
    rom_arr(integer(86)) <= "10011100101011011001100110001110";
    rom_arr(integer(85)) <= "01100110011010000111000001111000";
    rom_arr(integer(84)) <= "01110001011100110110100101100111";
    rom_arr(integer(83)) <= "01110010101001011001110010111011";
    rom_arr(integer(82)) <= "01111110100100001001110010010001";
    rom_arr(integer(81)) <= "10011101100001001001010110011100";
    rom_arr(integer(80)) <= "10010110101000011001011010110010";
    rom_arr(integer(79)) <= "10010111100001010111111101101110";
    rom_arr(integer(78)) <= "01100011011000000110110101110101";
    rom_arr(integer(77)) <= "01111000011101010111001001100111";
    rom_arr(integer(76)) <= "01110100011111010111100110000010";
    rom_arr(integer(75)) <= "10001110100001010111011001111110";
    rom_arr(integer(74)) <= "01101101011101110110011010000010";
    rom_arr(integer(73)) <= "01111101100000101000010110001000";
    rom_arr(integer(72)) <= "01110111101000000111011001101110";
    rom_arr(integer(71)) <= "01101000011011010110111101111000";
    rom_arr(integer(70)) <= "01110111011100110110111001110100";
    rom_arr(integer(69)) <= "01110100100001100110110010001000";
    rom_arr(integer(68)) <= "10000010100011011000101001111110";
    rom_arr(integer(67)) <= "10011011100010100111110001111111";
    rom_arr(integer(66)) <= "10000001100011100111111001111100";
    rom_arr(integer(65)) <= "01110101101001000111011101100110";
    rom_arr(integer(64)) <= "01100111011010100111001101110011";
    rom_arr(integer(63)) <= "01110011011100010110111101111001";
    rom_arr(integer(62)) <= "01111011011101111010110001101101";
    rom_arr(integer(61)) <= "01111111100011000111111010001110";
    rom_arr(integer(60)) <= "10000011100100001000010101100101";
    rom_arr(integer(59)) <= "01110111011110010111100010101000";
    rom_arr(integer(58)) <= "01100111011110010110111101100001";
    rom_arr(integer(57)) <= "01100100011100000111011101110111";
    rom_arr(integer(56)) <= "01110100011011010111000101101111";
    rom_arr(integer(55)) <= "01111100011101010111010110001111";
    rom_arr(integer(54)) <= "10000001100001101000101110011011";
    rom_arr(integer(53)) <= "10011011100011111001100110010011";
    rom_arr(integer(52)) <= "01111010011110100111100001110100";
    rom_arr(integer(51)) <= "01101111011100000101101001100100";
    rom_arr(integer(50)) <= "01101101011100100111000001110111";
    rom_arr(integer(49)) <= "01110101011100000111000001101101";
    rom_arr(integer(48)) <= "01101110011100010111011010010111";
    rom_arr(integer(47)) <= "01110111101000101001000110010111";
    rom_arr(integer(46)) <= "10001001100011111001101101111110";
    rom_arr(integer(45)) <= "10011010011100001001010101110100";
    rom_arr(integer(44)) <= "01101111011001110101111001101100";
    rom_arr(integer(43)) <= "01110101011100110111001001111001";
    rom_arr(integer(42)) <= "01110110011101010111001001101101";
    rom_arr(integer(41)) <= "01101001011001110111000001110100";
    rom_arr(integer(40)) <= "01110101011100100111001001101010";
    rom_arr(integer(39)) <= "10001001011001111000111010001111";
    rom_arr(integer(38)) <= "10111100011010010110111001101101";
    rom_arr(integer(37)) <= "01101011011100000111010001111001";
    rom_arr(integer(36)) <= "01110100011100110111010001110110";
    rom_arr(integer(35)) <= "01110111011101010111001101110010";
    rom_arr(integer(34)) <= "01110011011010110110011101101000";
    rom_arr(integer(33)) <= "01100100011011100110111101101111";
    rom_arr(integer(32)) <= "01110110011101000111000101101111";
    rom_arr(integer(31)) <= "01101110011011000110110001101110";
    rom_arr(integer(30)) <= "01110011011110000111010001110100";
    rom_arr(integer(29)) <= "01110100011100110111100101110100";
    rom_arr(integer(28)) <= "01110111011110010111011101110110";
    rom_arr(integer(27)) <= "01110001011101010111000101110010";
    rom_arr(integer(26)) <= "01110001011101000110111101101000";
    rom_arr(integer(25)) <= "01100110011010100110011101101010";
    rom_arr(integer(24)) <= "01101101011100100111001101110001";
    rom_arr(integer(23)) <= "01110010011110010111000101111001";
    rom_arr(integer(22)) <= "01110100011101110111011101110111";
    rom_arr(integer(21)) <= "01110111011101110111011001110100";
    rom_arr(integer(20)) <= "01110001011101000111001001110100";
    rom_arr(integer(19)) <= "01110101011101010111001001110010";
    rom_arr(integer(18)) <= "01110011011101010111000101110101";
    rom_arr(integer(17)) <= "01110100011100010111001001110101";
    rom_arr(integer(16)) <= "01110011011100100111100001111001";
    rom_arr(integer(15)) <= "01111001011110000111100001111000";
    rom_arr(integer(14)) <= "01110101011110010111011001110111";
    rom_arr(integer(13)) <= "01110101011101010111011101110010";
    rom_arr(integer(12)) <= "01110100011101010111100001110000";
    rom_arr(integer(11)) <= "01110101011110000111100001110010";
    rom_arr(integer(10)) <= "01110001011100110111010101110011";
    rom_arr(integer(9)) <= "01110010011101010111100001110110";
    rom_arr(integer(8)) <= "01110100011100010111001001110010";
    rom_arr(integer(7)) <= "01110101011101110111000101110100";
    rom_arr(integer(6)) <= "01110100011100100111010101110111";
    rom_arr(integer(5)) <= "01111001011110100111100001110011";
    rom_arr(integer(4)) <= "01111001011100110111100101110001";
    rom_arr(integer(3)) <= "01110010011100100111011101110110";
    rom_arr(integer(2)) <= "01110101011101000111011101110100";
    rom_arr(integer(1)) <= "01110010011110010111010101110110";
    rom_arr(integer(0)) <= "01100011000000000000000000000000";

    -- here ends the generated array allocation

    out_weights <= rom_arr(to_integer(unsigned(rom_index)));
end RTL;
