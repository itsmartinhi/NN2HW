library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
    port (
        in_rom_input_index:     in std_logic_vector(7 downto 0); -- the given rom input index
        in_rom_neuron_index:    in std_logic_vector(3 downto 0); -- the given neuron index
        out_data_rom:           out std_logic_vector(31 downto 0) -- the output datastream
    );
end ROM;

architecture RTL of ROM is 
    type t_rom_arr is array (0 to 2500) of std_logic_vector (31 downto 0);
    constant rom_arr: t_rom_arr := (
        -- here follows the generated array allocation
		2500 => "01110101011110000111100101110111",
		2499 => "01111000011101100111100001111000",
		2498 => "01110000011101000111001001110001",
		2497 => "01111011011101100110100101111010",
		2496 => "01110011011101110111011101111000",
		2495 => "01111001011101100111001101111000",
		2494 => "01110011011110100111100001110110",
		2493 => "01111001011101010111010001110111",
		2492 => "01111010011101111000100010001101",
		2491 => "10001101101001001001011010011100",
		2490 => "10010111101110001010010010101111",
		2489 => "10100001101001011010110010100010",
		2488 => "10100001100110101000111001111110",
		2487 => "01110111011100110111001001110110",
		2486 => "01110011011101000111011001101110",
		2485 => "01111011011101101001001010011100",
		2484 => "10001101100100101001010110011101",
		2483 => "10010011101010101001100110100101",
		2482 => "10100000101001011001001010011101",
		2481 => "10010000100100001001110001110111",
		2480 => "01110001011100010111011001111000",
		2479 => "01110010011100100111000001101011",
		2478 => "10001011100011111000011110001111",
		2477 => "10001001100010001000101010000110",
		2476 => "10000001011001110111000101110010",
		2475 => "10000000100010110110101110010001",
		2474 => "10000011011111000111100101110111",
		2473 => "01110001011110010111011101110010",
		2472 => "01110100011100010111010010000101",
		2471 => "10000110100111001000101001111100",
		2470 => "01111110011110000111001001110011",
		2469 => "01101101011111110111000101101111",
		2468 => "01110000011100100110100010000001",
		2467 => "01101111011011000110100101100111",
		2466 => "01110001011101000111000001110010",
		2465 => "01110110011101100111011110000000",
		2464 => "10000101011100100110110101111000",
		2463 => "01101000011011110110111001101100",
		2462 => "01011101011110010110100001111001",
		2461 => "01110110100001110110111110001011",
		2460 => "01110100011100100110011001101110",
		2459 => "01110110011101100111101001111001",
		2458 => "01110101011100110111010010000100",
		2457 => "01110101011010000111011101110100",
		2456 => "01110100011010110110100001110000",
		2455 => "01100100010111000101111001100011",
		2454 => "01100011011011010111000101110001",
		2453 => "01110100011111100111100001101110",
		2452 => "01101110011101110111000101110001",
		2451 => "01111001011101110111101010000100",
		2450 => "01110100011011110110100001110000",
		2449 => "01111001011100010111100001110111",
		2448 => "01100100011011000110101101011001",
		2447 => "01011011011001110110110001110010",
		2446 => "01101111011101010111111101101101",
		2445 => "01100101011100100111000101110001",
		2444 => "01110011011101000110110101101101",
		2443 => "01100111011010010111000001111110",
		2442 => "10000010011101000110011101110101",
		2441 => "01100100011010000110110001110101",
		2440 => "01101000011011100110111001111001",
		2439 => "10001010011111010110100101100011",
		2438 => "01101000011101000111001001110101",
		2437 => "01110011011100010110110101010110",
		2436 => "01011011011011010111010010000011",
		2435 => "01101111011100100111111101111011",
		2434 => "01111110100011010110101001101000",
		2433 => "10010100101010010111000001110001",
		2432 => "01111101100010010110011101100011",
		2431 => "01101000011101000111011101110100",
		2430 => "01110101011101100110110101011001",
		2429 => "01100001011011110111010001110100",
		2428 => "01110001011111101000000101111011",
		2427 => "10010000011101111000010010000111",
		2426 => "01110000100011000111100110010001",
		2425 => "10001011011100000111000001100100",
		2424 => "01101010011100100111100101110101",
		2423 => "01111010011100110110010001010110",
		2422 => "01100001100001000111000101111001",
		2421 => "01101011100000111000111110001011",
		2420 => "01111010011111000111001101110111",
		2419 => "10001011100001110111000110001111",
		2418 => "01111100011101001000001110000001",
		2417 => "01110000011100000111001101110010",
		2416 => "01110100011011100110110001010100",
		2415 => "01100110011110110111000110000100",
		2414 => "10001100100000001001110110001100",
		2413 => "10001101011011100111101101110100",
		2412 => "10001001100000110111101010001000",
		2411 => "10000010100001000111111010000011",
		2410 => "01110100011011000111100101111000",
		2409 => "01110111011100010110100101010001",
		2408 => "01011110011111101001010010010001",
		2407 => "01111111100001101001010010001111",
		2406 => "10001010011111001000111010000001",
		2405 => "10000000100000110111110101110101",
		2404 => "10000010101000010111111110010010",
		2403 => "01110100011100000111011001110100",
		2402 => "01110110011011000110000001010011",
		2401 => "01101010100001111001110010011000",
		2400 => "10011110100010001000101010011110",
		2399 => "10010001100010011000111101111001",
		2398 => "10000101100001000111100010001111",
		2397 => "10100000011111111001001010110011",
		2396 => "01101110011001110111001001111001",
		2395 => "01110111011011110110101001100000",
		2394 => "10100110101001101010101010001000",
		2393 => "10010101100101011000110010001110",
		2392 => "10010111100011001000010001110101",
		2391 => "10010111100100111001011110010111",
		2390 => "10011100101011011001100110001110",
		2389 => "01100110011010000111000001111000",
		2388 => "01110001011100110110100101100111",
		2387 => "01110010101001011001110010111011",
		2386 => "01111110100100001001110010010001",
		2385 => "10011101100001001001010110011100",
		2384 => "10010110101000011001011010110010",
		2383 => "10010111100001010111111101101110",
		2382 => "01100011011000000110110101110101",
		2381 => "01111000011101010111001001100111",
		2380 => "01110100011111010111100110000010",
		2379 => "10001110100001010111011001111110",
		2378 => "01101101011101110110011010000010",
		2377 => "01111101100000101000010110001000",
		2376 => "01110111101000000111011001101110",
		2375 => "01101000011011010110111101111000",
		2374 => "01110111011100110110111001110100",
		2373 => "01110100100001100110110010001000",
		2372 => "10000010100011011000101001111110",
		2371 => "10011011100010100111110001111111",
		2370 => "10000001100011100111111001111100",
		2369 => "01110101101001000111011101100110",
		2368 => "01100111011010100111001101110011",
		2367 => "01110011011100010110111101111001",
		2366 => "01111011011101111010110001101101",
		2365 => "01111111100011000111111010001110",
		2364 => "10000011100100001000010101100101",
		2363 => "01110111011110010111100010101000",
		2362 => "01100111011110010110111101100001",
		2361 => "01100100011100000111011101110111",
		2360 => "01110100011011010111000101101111",
		2359 => "01111100011101010111010110001111",
		2358 => "10000001100001101000101110011011",
		2357 => "10011011100011111001100110010011",
		2356 => "01111010011110100111100001110100",
		2355 => "01101111011100000101101001100100",
		2354 => "01101101011100100111000001110111",
		2353 => "01110101011100000111000001101101",
		2352 => "01101110011100010111011010010111",
		2351 => "01110111101000101001000110010111",
		2350 => "10001001100011111001101101111110",
		2349 => "10011010011100001001010101110100",
		2348 => "01101111011001110101111001101100",
		2347 => "01110101011100110111001001111001",
		2346 => "01110110011101010111001001101101",
		2345 => "01101001011001110111000001110100",
		2344 => "01110101011100100111001001101010",
		2343 => "10001001011001111000111010001111",
		2342 => "10111100011010010110111001101101",
		2341 => "01101011011100000111010001111001",
		2340 => "01110100011100110111010001110110",
		2339 => "01110111011101010111001101110010",
		2338 => "01110011011010110110011101101000",
		2337 => "01100100011011100110111101101111",
		2336 => "01110110011101000111000101101111",
		2335 => "01101110011011000110110001101110",
		2334 => "01110011011110000111010001110100",
		2333 => "01110100011100110111100101110100",
		2332 => "01110111011110010111011101110110",
		2331 => "01110001011101010111000101110010",
		2330 => "01110001011101000110111101101000",
		2329 => "01100110011010100110011101101010",
		2328 => "01101101011100100111001101110001",
		2327 => "01110010011110010111000101111001",
		2326 => "01110100011101110111011101110111",
		2325 => "01110111011101110111011001110100",
		2324 => "01110001011101000111001001110100",
		2323 => "01110101011101010111001001110010",
		2322 => "01110011011101010111000101110101",
		2321 => "01110100011100010111001001110101",
		2320 => "01110011011100100111100001111001",
		2319 => "01111001011110000111100001111000",
		2318 => "01110101011110010111011001110111",
		2317 => "01110101011101010111011101110010",
		2316 => "01110100011101010111100001110000",
		2315 => "01110101011110000111100001110010",
		2314 => "01110001011100110111010101110011",
		2313 => "01110010011101010111100001110110",
		2312 => "01110100011100010111001001110010",
		2311 => "01110101011101110111000101110100",
		2310 => "01110100011100100111010101110111",
		2309 => "01111001011110100111100001110011",
		2308 => "01111001011100110111100101110001",
		2307 => "01110010011100100111011101110110",
		2306 => "01110101011101000111011101110100",
		2305 => "01110010011110010111010101110110",
		2304 => "01100011000000000000000000000000",
		2244 => "01111001011110010111100001110111",
		2243 => "01110011011101100111000101110011",
		2242 => "01110101011110010111001101110101",
		2241 => "01110001011101100111100101110101",
		2240 => "01111001011101010111100001110100",
		2239 => "01111010011101110111010001110011",
		2238 => "01110010011110000111101001110011",
		2237 => "01110110011101100111010001110110",
		2236 => "01110001011101000111000001101010",
		2235 => "01101111011100010111000101101010",
		2234 => "01100111011010110111010001110100",
		2233 => "01110011011011000111000101110100",
		2232 => "01110101011010110111010101110111",
		2231 => "01110110011101110111100001110011",
		2230 => "01110100011101100111100101110100",
		2229 => "01101101011100110110111101111011",
		2228 => "10001001100001011010101110100000",
		2227 => "10100110101001100111110010001101",
		2226 => "10101011101001000111000101110000",
		2225 => "01110001011100000110001001101101",
		2224 => "01111001011100110111100101110011",
		2223 => "01110001011100100111010101101100",
		2222 => "01110001011100000111001010001000",
		2221 => "10111111100111100110011111001000",
		2220 => "10001010101010001001001010010101",
		2219 => "10100011011111011000001110011111",
		2218 => "01110000011001100101110001100110",
		2217 => "01101011011101100111011101110110",
		2216 => "01110101011101010111001001101110",
		2215 => "10000100100000001000000110001000",
		2214 => "10010101101000010111101010000110",
		2213 => "10000101011110111001011110000101",
		2212 => "10000010011111000111111010011111",
		2211 => "01101011011010000110101101110100",
		2210 => "01110100011110010111011001111001",
		2209 => "01110111011100100111000001101110",
		2208 => "01111101011110111000101001101011",
		2207 => "01110100011111110111110001110100",
		2206 => "01111111100001010111100101111101",
		2205 => "10000011011110100111100001101110",
		2204 => "10001010100011010111100001111101",
		2203 => "01110101011100010111001101110001",
		2202 => "01110100011101100110111101100010",
		2201 => "01110110100011110110111110001110",
		2200 => "01111111011111101001000101110010",
		2199 => "01110011011101111000001001101000",
		2198 => "01111101011010111001010101110110",
		2197 => "10100011101000000111010001110110",
		2196 => "01101010011101100111011001110101",
		2195 => "01110111011101100110100101100111",
		2194 => "10001010100011001011000110011101",
		2193 => "10001010011110000111100101101010",
		2192 => "10000010011001011000001001111110",
		2191 => "01110101100100100111110010001000",
		2190 => "10101001011110010111011001101111",
		2189 => "01100110011100010111001101111000",
		2188 => "01110110011100100110010001101011",
		2187 => "10100110101000100110101101110100",
		2186 => "10000000100010001000001101111110",
		2185 => "01110010011100100111001110000011",
		2184 => "01110011100011101000111010000011",
		2183 => "01101111100001101010010001101110",
		2182 => "01100111011101000111001101110010",
		2181 => "01111001011101000110001001110001",
		2180 => "10010000011100110110111110000011",
		2179 => "01110001011101100110110101110011",
		2178 => "01110110011101011000010110001101",
		2177 => "10010111100101101001001101111111",
		2176 => "01110100100110000111010001101100",
		2175 => "01101100011101000111010101110011",
		2174 => "01111000011100000110001010000111",
		2173 => "10001110011101010111101101110101",
		2172 => "01110111011001100111011110000110",
		2171 => "01110000100000111000100110010001",
		2170 => "10001100100000111001110110001011",
		2169 => "10110011011100000111000101110010",
		2168 => "01110101011101100111010101110011",
		2167 => "01110100011011110110100001101010",
		2166 => "10000100011011000111000101101101",
		2165 => "01100111011100111000100010001000",
		2164 => "01111110100001101000101010011001",
		2163 => "10000101100100100111110101110101",
		2162 => "01110100011101010110101101101000",
		2161 => "01111010011101010111001001110110",
		2160 => "01110110011100000111101001100101",
		2159 => "01101010011101000111001101110000",
		2158 => "01111001100001000111011101111001",
		2157 => "10000001100110101001000010001101",
		2156 => "01111001011101011000011001110001",
		2155 => "01110101011100110110011101101001",
		2154 => "01110011011101100111010101111001",
		2153 => "01110011011101010111101101100111",
		2152 => "01100011011001110111010001101011",
		2151 => "01111101011101001000001110000010",
		2150 => "10000011100010101001100110001110",
		2149 => "10011100100000010110100101101011",
		2148 => "01101101011110010111100001100101",
		2147 => "01110111011101000111011101110000",
		2146 => "01111000011101010111110110010000",
		2145 => "10011100100010000110101010101100",
		2144 => "01110110011111010110111110001000",
		2143 => "10011001011101111010100010011001",
		2142 => "10010000011011101000000001111110",
		2141 => "01111011100110001000001001110010",
		2140 => "01111011011101110111100101110000",
		2139 => "01110000011101110111100110111100",
		2138 => "10110001101000011011000110001001",
		2137 => "10011100011100111000011101111101",
		2136 => "10000111100001101001111010001101",
		2135 => "10000111011111001000110001101101",
		2134 => "10100100011100001010010001111000",
		2133 => "01111110011110010111011101110100",
		2132 => "01110101100001100111100110010111",
		2131 => "10010110100100010111100110000000",
		2130 => "01110101011010010111000001111001",
		2129 => "01111110101101001001101010001111",
		2128 => "10001011100100101010001010100110",
		2127 => "11000110100010101000111010000001",
		2126 => "01110001011100010111011001110101",
		2125 => "01110101011110100111001001110110",
		2124 => "10010011100100001001001110010000",
		2123 => "10011101100100110111011001101100",
		2122 => "01011110011101010111100110011011",
		2121 => "10000011100110001000100101111010",
		2120 => "01110101100001000111010010010010",
		2119 => "01101110011100110111011001110100",
		2118 => "01110010100100001001011110011100",
		2117 => "10011010100010011000111010000001",
		2116 => "10000001011101101000101101111100",
		2115 => "01100101011101110111110001101001",
		2114 => "10000111011110001000101110010000",
		2113 => "01111110100100110111011101110110",
		2112 => "01110010011101100111010001110110",
		2111 => "01111111100010011001000110110011",
		2110 => "10001010100001011000111110000010",
		2109 => "10010010100010110111011110001111",
		2108 => "01110011011011101000101110000110",
		2107 => "01111001100010101000101101110001",
		2106 => "10011011100101101000100101111001",
		2105 => "01111100011100110111010001110001",
		2104 => "01110011011101100111111010011001",
		2103 => "10101000011111001001010001110010",
		2102 => "01110111100010000110111001111011",
		2101 => "10001110011000000111110101101110",
		2100 => "01101101100001000111001110100111",
		2099 => "01101100011011100111010101110010",
		2098 => "01110000011100010111011101110001",
		2097 => "01110010011101111001001101110001",
		2096 => "10011101011101010111011110000001",
		2095 => "10011111011011111000110101111110",
		2094 => "10001111100000001000000010011011",
		2093 => "01110101011110101000001001111010",
		2092 => "01110011011011110110111001101111",
		2091 => "01110110011100100111011001110100",
		2090 => "01111000011101101000111010000011",
		2089 => "01101101011101110111111010010111",
		2088 => "10001000011011011010000010000111",
		2087 => "01111111100010011000000010010000",
		2086 => "10100011011011011000011001110001",
		2085 => "10000010011011000110101101110101",
		2084 => "01110000011101100111100001110110",
		2083 => "01111000011111001000010110000110",
		2082 => "01111110100100001000000110100111",
		2081 => "01110010101110011000101110110011",
		2080 => "10100001110001010110010011011101",
		2079 => "10001011100111001001000010000101",
		2078 => "01110010011011000111000101110011",
		2077 => "01110110011100100111010101110100",
		2076 => "01111000011100010111010001110101",
		2075 => "10000010100010000111110101110010",
		2074 => "01110001100011101000001101110110",
		2073 => "01110110011101010111100101110011",
		2072 => "01110100011110010111010101111000",
		2071 => "01110001011100100111001001110001",
		2070 => "01110010011101010111100101110110",
		2069 => "01110011011101000111001001111001",
		2068 => "01110101011100110111001001110101",
		2067 => "01110011011101010110111001101110",
		2066 => "01110000011100110111000101110000",
		2065 => "01110000011100000111100001110100",
		2064 => "01110011011110010111000101110110",
		2063 => "01110110011100100111010101110010",
		2062 => "01110011011101110111010001111001",
		2061 => "01110100011100010111011101110011",
		2060 => "01111000011100010111010101110110",
		2059 => "01110110011101110111100001110011",
		2058 => "01110010011101000111100101111000",
		2057 => "01111010011100100111100101110001",
		2056 => "01111001011100100111011101111000",
		2055 => "01110001011100100111001001110011",
		2054 => "01110010011101000111011001111010",
		2053 => "01110001011101010111100101111000",
		2052 => "01110111011101000111011101110101",
		2051 => "01110110011100000111001001110100",
		2050 => "01110011011101000111001001111001",
		2049 => "01111000011101100111000101110001",
		2048 => "00000000000000000000000000000000",
		1988 => "01111001011100110111001101110110",
		1987 => "01110100100000001000000001111011",
		1986 => "10000011100001001000000101111111",
		1985 => "01111100100000011000011001111011",
		1984 => "01111001011111000111010101111000",
		1983 => "01110011011101110111000101110010",
		1982 => "01110111011110100111011001110011",
		1981 => "01110001011110010111011001110000",
		1980 => "01110100100000100111100001110110",
		1979 => "10010110100101101001011110001100",
		1978 => "10011101100101011001010110000001",
		1977 => "10000101100011011000110010000100",
		1976 => "01111011011000100110100001101111",
		1975 => "01111001011110000111100101110110",
		1974 => "01110001011110000111011101110001",
		1973 => "01110001011101010111010101110000",
		1972 => "01111111100100011001000010011000",
		1971 => "10011010101000001001100010101110",
		1970 => "10110110100101111010000110010100",
		1969 => "10000100011100110111011010000100",
		1968 => "01110111011101010111010001110111",
		1967 => "01110100011101100110111101101110",
		1966 => "01011011011001010110100001101011",
		1965 => "01101101011010001000010101110011",
		1964 => "01111001011110111000111101110000",
		1963 => "01111101100000010111010110001011",
		1962 => "10001110100101111001101101111111",
		1961 => "01110111011101010111001101110101",
		1960 => "01110001011100010111010001101111",
		1959 => "01010110010101000101000101011001",
		1958 => "01101000011011010111001001110000",
		1957 => "01111010011011100110001001100100",
		1956 => "01100111011011100110111001011101",
		1955 => "10011100100011110111101001110010",
		1954 => "01100011011100110111011001111001",
		1953 => "01110001011100110111010101101111",
		1952 => "01011001010100010101011101100011",
		1951 => "01110101011010110110101001110111",
		1950 => "01110000011101110110000001111101",
		1949 => "01100111011101010111001001110111",
		1948 => "10000001011100010111000101011110",
		1947 => "01100010011010010111010101111010",
		1946 => "01110110011100110111000001110100",
		1945 => "01010111010100000101101001100101",
		1944 => "01100110011010000110100101110100",
		1943 => "01101000010111110110010001110001",
		1942 => "01101111011101010110111101110100",
		1941 => "01011101010111010110001101011010",
		1940 => "01101000011100000111010101110100",
		1939 => "01110100011101010110110001101110",
		1938 => "01100010010100010101111001011010",
		1937 => "01100111010110100110000101100000",
		1936 => "01100110011110110111010001111011",
		1935 => "01101110011011100110111001110011",
		1934 => "01100110010110110110001001011110",
		1933 => "01100110011100010111010001110001",
		1932 => "01110111011110010111010101101111",
		1931 => "01010101010110100110111001110001",
		1930 => "01110010011001000110101001101000",
		1929 => "01101000011111100110111001110100",
		1928 => "01110001011000000111001101110011",
		1927 => "01100111011011000110111101110100",
		1926 => "01101101011111000111011001110110",
		1925 => "01111001011101010111011101101101",
		1924 => "01011101011101011000000001110011",
		1923 => "01110100011101100111011101110010",
		1922 => "01110001011100101000001101101110",
		1921 => "01111000011101000110111101101110",
		1920 => "01101100011001110111111101111101",
		1919 => "01101110011101110111010001110001",
		1918 => "01110000011101110111110110000010",
		1917 => "01110110100000000111010110001100",
		1916 => "01101110100011010111011001110111",
		1915 => "10001000100001011000000110000110",
		1914 => "01101101011001110111001001110100",
		1913 => "01101111011101011000000010000010",
		1912 => "01101010011100010111011001110001",
		1911 => "01110001011011110110011101101000",
		1910 => "01110010011100101001010110011000",
		1909 => "10010010011110111001100001111000",
		1908 => "10001011010110010111110101101110",
		1907 => "01011010011010000111000001111001",
		1906 => "10100111011101110110111001111101",
		1905 => "01101101011101110111001101110100",
		1904 => "01110010011011100110000001101011",
		1903 => "10010111101000011000111110010110",
		1902 => "01111011101000111100000001011111",
		1901 => "10001100011001100110110001011100",
		1900 => "01100111011100010110101101101100",
		1899 => "01110001011110100111001101110000",
		1898 => "10000011011101110111000001110110",
		1897 => "01110010011110000110111001110010",
		1896 => "10010100100010100111000110011111",
		1895 => "11000011100011011000100110001001",
		1894 => "01110001011100010110001001011001",
		1893 => "01100011011101000111000101111010",
		1892 => "01110110011101101001000110001001",
		1891 => "10001001100000000111101001110100",
		1890 => "01110011011101010111110001111010",
		1889 => "01101100011110011010000010010000",
		1888 => "01100111011100110111101010001110",
		1887 => "01111010011100010101100101001111",
		1886 => "01110000100001100111000001101000",
		1885 => "10000000101100101000001110001110",
		1884 => "10011000100010100111011001111000",
		1883 => "01110011011111010111011001100101",
		1882 => "01101110101010111000111001111001",
		1881 => "01111010101000001001011110100111",
		1880 => "10101011011011010101000001011101",
		1879 => "10011000011100010111000011011010",
		1878 => "10101001011110011000100010011110",
		1877 => "10100000100110010111111001110101",
		1876 => "01110111011100110110111001100101",
		1875 => "01110000100111001001001010101010",
		1874 => "10000010101010011000111110001011",
		1873 => "10100110101100111000100010000110",
		1872 => "10010100101101101001000001101110",
		1871 => "10010001100001100111111010001101",
		1870 => "10010001100110110111110001110101",
		1869 => "01110010011110110111011101101011",
		1868 => "01110111100111001001101010101011",
		1867 => "10100001100010111000011010110100",
		1866 => "10001100100010001001100001100111",
		1865 => "01100110011101101001000101111000",
		1864 => "10000110100011101000110110001111",
		1863 => "10010001100010110111111101110010",
		1862 => "10000000011101010111100001111100",
		1861 => "10000011100100011001011101110110",
		1860 => "10010100100101111011010110001111",
		1859 => "10010100101010010111100110100011",
		1858 => "10000010011110001000110010000111",
		1857 => "10000110100100111000101010010001",
		1856 => "10001111100000000111110101110111",
		1855 => "01110101011101100110101001110010",
		1854 => "10001100100100100111010110010101",
		1853 => "10000010100111101000001010001000",
		1852 => "10011000100010100110111110011100",
		1851 => "10010010011111111001000110011000",
		1850 => "10100101100011101000101110001100",
		1849 => "10010101100000000111101001110010",
		1848 => "01110100011110010111001001111000",
		1847 => "10000000100000111000110110100100",
		1846 => "01110111101000111000101010001011",
		1845 => "10001001011011011000110110001111",
		1844 => "01111011100011101000110101111011",
		1843 => "10011001100011000111110110001010",
		1842 => "10010011011111110111010101111001",
		1841 => "01111000011110000111000101101101",
		1840 => "01100101011101001000011101110011",
		1839 => "01111001011111111000101010000101",
		1838 => "01111100011110110111010010010010",
		1837 => "10101110100011101000111010011010",
		1836 => "10010000100101011000110101111111",
		1835 => "10000110011101000111010001110101",
		1834 => "01110111011110000111000101110000",
		1833 => "01101111011010010110011101011011",
		1832 => "01100101011011100110111001110011",
		1831 => "01110001011100101000000110001011",
		1830 => "01110111011101101001010110010010",
		1829 => "10000100011110100111110001110010",
		1828 => "01110100011101000111100101110010",
		1827 => "01110101011101100111011101110001",
		1826 => "01110100011100010111010101101111",
		1825 => "01101010011010110110011101100110",
		1824 => "01100101011001010110100001100100",
		1823 => "01011100010101110101111101101001",
		1822 => "01101011011011000111010001110110",
		1821 => "01110001011100100111001101110101",
		1820 => "01110111011100110111100101110111",
		1819 => "01110111011110000111011001110111",
		1818 => "01110100011101110110111001110001",
		1817 => "01101101011011110110100101101011",
		1816 => "01101001011010000111001101110010",
		1815 => "01110101011101110111101001111000",
		1814 => "01110100011100010111001101111001",
		1813 => "01110011011101100111001101110101",
		1812 => "01110000011110010111001001110001",
		1811 => "01110010011101100111001001110101",
		1810 => "01110100011100010111010001110101",
		1809 => "01110100011100000111000001110111",
		1808 => "01110101011101110111010001111000",
		1807 => "01110101011101010111000101111000",
		1806 => "01110001011110010111100001110001",
		1805 => "01110001011100110111000101110111",
		1804 => "01110100011110010111011001110110",
		1803 => "01110100011110000111000101110100",
		1802 => "01110111011101110111101001111001",
		1801 => "01110001011101100111000101111001",
		1800 => "01111001011101110111100101110011",
		1799 => "01110011011110010111001001110110",
		1798 => "01110110011101000111000101110010",
		1797 => "01110000011101110111001001110001",
		1796 => "01110111011110000111011101110101",
		1795 => "01110100011100110111001001110001",
		1794 => "01110101011110010111000101110100",
		1793 => "01111001011101000111001101111001",
		1792 => "11010100000000000000000000000000",
		1732 => "01110111011110010111000101110011",
		1731 => "01110010011100100111010001110100",
		1730 => "01110011011101100111001101110011",
		1729 => "01111000011101000111010001111000",
		1728 => "01110111011101110111000101110101",
		1727 => "01110100011101110111100001111001",
		1726 => "01110110011100100111000101110010",
		1725 => "01110010011110000111000001110001",
		1724 => "01110001011101000111001001111001",
		1723 => "01110001011101100111100001111001",
		1722 => "01110011011101110111001101110010",
		1721 => "01111000011100010111010001110010",
		1720 => "01110010011101100111001101110010",
		1719 => "01111001011110010111010101110011",
		1718 => "01111000011100010111011001110000",
		1717 => "01110011011101010111100101110011",
		1716 => "01101111011100110111001101101111",
		1715 => "01101010011100000110110101110111",
		1714 => "01110101011100100111001101110101",
		1713 => "01110010011101110111000101110110",
		1712 => "01110110011100100111010101110010",
		1711 => "01110101011100100111100001110010",
		1710 => "01110010011100100111000101110000",
		1709 => "01101101011101010111100101111011",
		1708 => "01101111011010000110001101100101",
		1707 => "01011000011000000110010001101010",
		1706 => "01110010011101000111001101111001",
		1705 => "01110001011101000111100001110111",
		1704 => "01110001011110010111001001101101",
		1703 => "01101101011011100111011010000001",
		1702 => "10010010100101010111011101110100",
		1701 => "01110101011110110111010001110110",
		1700 => "01101111011010010111000001101010",
		1699 => "01100111011010110111001101110001",
		1698 => "01111000011101110111011101110000",
		1697 => "01111001011101100111100001100110",
		1696 => "01100100011010011000011110001100",
		1695 => "01111111011110110111011010000101",
		1694 => "10100111011010011001001010010001",
		1693 => "01101010100111101000011001111111",
		1692 => "01110101010111100110011101101011",
		1691 => "01110101011100110111100001110110",
		1690 => "01110111011101010110111001110000",
		1689 => "01101110100000110111001010010111",
		1688 => "10001111101000111001111110001000",
		1687 => "10001001100110111001010110100101",
		1686 => "10001100100011001000101110100111",
		1685 => "01111100011010100110011001101000",
		1684 => "01110101011100100111010101110101",
		1683 => "01110110011101000110110101101101",
		1682 => "10000000011110001001000110011010",
		1681 => "01111100100101001000001110001000",
		1680 => "10001110101000110111111110011111",
		1679 => "10010100101001101001111101101110",
		1678 => "10011101011101010111010001101110",
		1677 => "01110011011101010111100001110111",
		1676 => "01110011011100100110100001110011",
		1675 => "10001101100111001000100001111111",
		1674 => "10000101100001001000101110000011",
		1673 => "10001011100110011000011110100011",
		1672 => "10101010101000011001110001111000",
		1671 => "10001001100100010111100101110011",
		1670 => "01110010011110100111010101110110",
		1669 => "01110101011100101000001110000100",
		1668 => "10001001011101110111110101111010",
		1667 => "01111001100011001000101110001111",
		1666 => "01111001011101001001101010110000",
		1665 => "01111101100011111001000110001001",
		1664 => "10011110100000000111001001100000",
		1663 => "01110011011101100111001001110010",
		1662 => "01110101011010111000101010000110",
		1661 => "10000111100010111000010110000011",
		1660 => "10000110100000001000100001110101",
		1659 => "01110111100100001000100110000101",
		1658 => "10101100101011011001111110010110",
		1657 => "10001000100001011000001101011000",
		1656 => "01110000011101110111100001111000",
		1655 => "01101111011000111000100010000001",
		1654 => "01111000100001001000100101111011",
		1653 => "10001010100010100111001010000001",
		1652 => "01111101100010000111100001111001",
		1651 => "10110100100100011001110010001110",
		1650 => "10010110101001011000010101011011",
		1649 => "01101000011101010111011101110100",
		1648 => "01110111011000111000110010000110",
		1647 => "10000001011110111000110110000110",
		1646 => "01111010011110101000001001111011",
		1645 => "01111011100101111000101110010101",
		1644 => "10010001100010010111111110010001",
		1643 => "10010000100100000111000001011001",
		1642 => "01110001011110100111001001111000",
		1641 => "01110001011001100111111010010000",
		1640 => "10010001100011111000101001111001",
		1639 => "01111101011110000110010110001101",
		1638 => "01111111011100110111100110001011",
		1637 => "10100100100101101000111110001101",
		1636 => "01111010100100101000101001011110",
		1635 => "01110010011100010111011101110101",
		1634 => "01110010010110100101100110011001",
		1633 => "10110101100011101001011101111010",
		1632 => "10000100011100100110110001111101",
		1631 => "10000100011011111001011010010000",
		1630 => "01111001100011110111100101110110",
		1629 => "10001001101010011000100101110001",
		1628 => "01101111011101010111000101110010",
		1627 => "01110001010110000110000110011001",
		1626 => "10111101101001011001001001111001",
		1625 => "01100011011011010111010001111100",
		1624 => "01101010011011111001001010010001",
		1623 => "10100001100001111000111010010011",
		1622 => "10100010100011010111110001110011",
		1621 => "01101011011101100111011101110000",
		1620 => "01110100010110000101001001111000",
		1619 => "10011011011011101000010101111001",
		1618 => "01111010011001110110011101110101",
		1617 => "01011100011101001001011110010001",
		1616 => "01110111100000101001101110000110",
		1615 => "10010110011101000111110001110101",
		1614 => "01110010011100100111100101110100",
		1613 => "01110011011001100101100001110001",
		1612 => "01110100011001000111000101110010",
		1611 => "01101000011001010110011101100100",
		1610 => "01011100011001110111010001101101",
		1609 => "01101110011101110110111110000000",
		1608 => "01111111011100010110110001110010",
		1607 => "01101011011100110111001101110100",
		1606 => "01110000011001010101101101101000",
		1605 => "01101101011011010111101001101110",
		1604 => "01100100010110100101100101011101",
		1603 => "01100111011011110101110001101100",
		1602 => "01110000011001010110101101110000",
		1601 => "01111100011011100110100110000010",
		1600 => "01110100011100110111101001111001",
		1599 => "01101111011011000110010101100001",
		1598 => "01100101011011010111000101101010",
		1597 => "01100000010110100110110001101000",
		1596 => "01011100011000000111010001101001",
		1595 => "01101111011100000111100001110010",
		1594 => "01110000011011100111010001110111",
		1593 => "01101101011101010111010101110101",
		1592 => "01110101011100110111000010001000",
		1591 => "01110101011011100111010001101001",
		1590 => "01101000011010000110101101100111",
		1589 => "01110001011100110110001101110001",
		1588 => "01111010011100000111010101110011",
		1587 => "01111111011000100111011001110011",
		1586 => "01101111011110000111000101111001",
		1585 => "01110110011110110111010110001110",
		1584 => "10001000011100100111010101101111",
		1583 => "01101000011001100110111101101010",
		1582 => "01110110011010000110011101110000",
		1581 => "01101110011010000111010101110111",
		1580 => "01110101011000110110110001110101",
		1579 => "01101111011110000111010001111000",
		1578 => "01111010011101110111001001111111",
		1577 => "10011110011100101000101010000110",
		1576 => "10011010100011011000010001110011",
		1575 => "01101101100000010110110001110101",
		1574 => "01101011100011110111101110000110",
		1573 => "01101100011100100110100001110110",
		1572 => "01101111011100100111010101110110",
		1571 => "01111010011110000110101101100000",
		1570 => "10001011100011001000011110000101",
		1569 => "10000000100000011001000110010011",
		1568 => "10000010100001011000001101111111",
		1567 => "01111101100001110111000110000001",
		1566 => "01110101011111010111100001111011",
		1565 => "01110100011110010111001001110111",
		1564 => "01110011011101010110110010000001",
		1563 => "10001101100001100111111101111001",
		1562 => "10001101100010000111110110000011",
		1561 => "10001100100011001001000010001100",
		1560 => "10010000100011111001000110001000",
		1559 => "10000111100000010111010001110110",
		1558 => "01111000011100110111010001110010",
		1557 => "01110111011110000111000101110110",
		1556 => "01111110100001101000111110000111",
		1555 => "10001100100001001000010110000011",
		1554 => "10000011100010111000101010010011",
		1553 => "10010100100100111000100110001111",
		1552 => "10001100011111100111001001111010",
		1551 => "01110111011100000111000001111001",
		1550 => "01110111011100100111001001111001",
		1549 => "01111100011110100111101001111000",
		1548 => "01111110011111000111011101110101",
		1547 => "01111000011110001000001010000111",
		1546 => "01111011011110100111110010000000",
		1545 => "01111111011111010111100001111001",
		1544 => "01110001011110010111001101111000",
		1543 => "01110111011101010111001001110100",
		1542 => "01111001011110010111000101110110",
		1541 => "01110100011110010111010101110110",
		1540 => "01110011011100110111001001111001",
		1539 => "01110101011100010111000001110110",
		1538 => "01110010011100100111011001110101",
		1537 => "01110011011101000111001001110101",
		1536 => "01101111000000000000000000000000",
		1476 => "01110010011100010111010101110010",
		1475 => "01110011011101100111011101110100",
		1474 => "01110100011101010111011101110010",
		1473 => "01110010011100110111000101111001",
		1472 => "01110010011101100111000101110010",
		1471 => "01110110011101000111010001110001",
		1470 => "01110110011110010111001101110111",
		1469 => "01110101011101010111001001110111",
		1468 => "01110111011100110111011101111010",
		1467 => "01110010011010010111000001111011",
		1466 => "10001011011111010111111110001100",
		1465 => "10000001011101010110100001100101",
		1464 => "01100111011011010111011001110110",
		1463 => "01110111011110010111011101110101",
		1462 => "01110001011101000111011110000001",
		1461 => "10001011100011011000111010000001",
		1460 => "10001100100101011010000110101111",
		1459 => "10111000011111111011000110101010",
		1458 => "10101011100111101001111001111000",
		1457 => "01111001011111010111010110000001",
		1456 => "01111001011110010111011001110101",
		1455 => "01110100011110100111000101111010",
		1454 => "01111111100010110111011010001001",
		1453 => "10000001101000101010110110000000",
		1452 => "10100001101000011010011110001101",
		1451 => "10001011100001111010011110001010",
		1450 => "01111011011111000111110101111011",
		1449 => "01111001011101010111011001110100",
		1448 => "01110011011101000111100010000000",
		1447 => "10000101100000000111100110001101",
		1446 => "01110111011011110111011110001011",
		1445 => "01110010100000110111001010000110",
		1444 => "10000001101001000111011110011001",
		1443 => "01101101100001111001000010000111",
		1442 => "01111111011110000111011101111000",
		1441 => "01110110011101001000000010001011",
		1440 => "10010010100010110111101110000101",
		1439 => "10001101100110100111011110000111",
		1438 => "01111110100010001000000010000000",
		1437 => "01111110011100010111111101111011",
		1436 => "10000011011100010110110110010100",
		1435 => "01111010011100100111100001111001",
		1434 => "01110100011101000111110010000100",
		1433 => "10000111100110111001101010011110",
		1432 => "01111110100000001000110001110010",
		1431 => "01111110100000100111101001111100",
		1430 => "10001011011111101000010010001001",
		1429 => "10100100100100100111101110010000",
		1428 => "01111001011100000111001101110100",
		1427 => "01111001011100111000000001111100",
		1426 => "10000111101011000111110001111111",
		1425 => "10010110100010011000111110001011",
		1424 => "01110101011100111000100001111000",
		1423 => "10001010100000001010000110010110",
		1422 => "01111000100100011010011101111111",
		1421 => "10000010100000000111010101111000",
		1420 => "01110100011100010111000110001001",
		1419 => "10010101100000101001001010011100",
		1418 => "01110011100010000111001001110000",
		1417 => "01111101011011101000100110000000",
		1416 => "10000110100011100111010010101000",
		1415 => "01110110100110100111010010100101",
		1414 => "01111100011111100111010101110110",
		1413 => "01110110011011110110100110001110",
		1412 => "10010000100011000111011101110001",
		1411 => "10000001011010011000100101111111",
		1410 => "01111111011111110111100101110011",
		1409 => "01111110011110110111010101110101",
		1408 => "10010010101101101001000110100111",
		1407 => "01111011011101110111100001111001",
		1406 => "01110101011100000110010001111010",
		1405 => "10001100011100001000010001111111",
		1404 => "01111111100110101001000101111111",
		1403 => "01111000011010010110100001100111",
		1402 => "01110001011101010111011101110100",
		1401 => "01101101101001111000100101111101",
		1400 => "01111010011010110111001001111001",
		1399 => "01110000011010110110101101111101",
		1398 => "10001111101001010111100110011001",
		1397 => "10000000011001100111100101101000",
		1396 => "01111010011011110111101101111011",
		1395 => "01110110100000000110100001110000",
		1394 => "01101000011011110111001001101111",
		1393 => "01110100011100110111011101110101",
		1392 => "01101110011011010110011010010010",
		1391 => "10001101011001011000100101110111",
		1390 => "01111001100111010111000101111010",
		1389 => "01101101011011100111110010001110",
		1388 => "10000010100001111000111001111001",
		1387 => "01101111011110110110111101110011",
		1386 => "01101111011100110111100101111000",
		1385 => "01110100011100100101100101110111",
		1384 => "01110100100010100111000101111100",
		1383 => "01100111011010010110100101110000",
		1382 => "01110111011111010111111010001010",
		1381 => "10000001100110011000000010000000",
		1380 => "10000001011101010111001110000000",
		1379 => "01110101011101010111001001110111",
		1378 => "01110011011100110101111100111000",
		1377 => "01011001011011010110111110000111",
		1376 => "10000011011100110111001001100101",
		1375 => "01101011011101111001101010101000",
		1374 => "10010110100000010111111101111010",
		1373 => "10100001011100101001011110000100",
		1372 => "01110010011101000111010101110001",
		1371 => "01110101100011000111010100101011",
		1370 => "00111110010101000101111101101111",
		1369 => "01100111011010010110010001101100",
		1368 => "10001000011101001001011110001111",
		1367 => "10001110101000010111110110000100",
		1366 => "10001110101001010111010101110111",
		1365 => "01101100011101110111011101110100",
		1364 => "01110001100010111101001011000101",
		1363 => "01110011010111000110100001100111",
		1362 => "01101001011100100110111101110100",
		1361 => "01110010100001101010111010001011",
		1360 => "10001011100001001000100110010010",
		1359 => "10010000100101100111011001110100",
		1358 => "01100010011101000111100101111010",
		1357 => "01111010100101011110000011110011",
		1356 => "10111110011010010111001001110000",
		1355 => "01101111011010100110100001101101",
		1354 => "01110100011110101000011010011000",
		1353 => "10000110100101011010000110011100",
		1352 => "10010100011011100111001001110000",
		1351 => "01100111011101000111011101111000",
		1350 => "01110111100010111011101111010111",
		1349 => "10011000100111111011011001110101",
		1348 => "01110101100000110111100101100111",
		1347 => "01100110011100000111001001111111",
		1346 => "10010001011111100110110001111100",
		1345 => "01110100100000010110111001010100",
		1344 => "01100010011100000111001001110011",
		1343 => "01110101100010001011001111000110",
		1342 => "10110001011100111000100010010111",
		1341 => "10001100011110011000000001111110",
		1340 => "01110000011100110111001101111000",
		1339 => "10000000100000111000100101111110",
		1338 => "01101101011110100110101001000010",
		1337 => "01100101011110000111000101110111",
		1336 => "01111000011111101010110010101011",
		1335 => "10010111100101011000100001111110",
		1334 => "01110101100000110111110110000011",
		1333 => "01100100100001110110101010000010",
		1332 => "01111101100101100111010010110001",
		1331 => "01111001011111000110110001001110",
		1330 => "01101000011101010111100101110110",
		1329 => "01110110100001001001011110100101",
		1328 => "10001011100011110111000110001001",
		1327 => "10011010100000010111110101110111",
		1326 => "01111000100010110111100010000101",
		1325 => "01111000011101100111011001111001",
		1324 => "01110111011101010111001001100000",
		1323 => "01100110011110010111100101111000",
		1322 => "01110010011111011001001010010100",
		1321 => "10001100100011100111101010100100",
		1320 => "01110100100001011001000110000011",
		1319 => "01101100011101011000001001111111",
		1318 => "10001000100111110111011001110011",
		1317 => "01110100011000100110001001011111",
		1316 => "01101111011101000111011001111001",
		1315 => "01110011011110001000101110011100",
		1314 => "10001110100000011001011101101011",
		1313 => "10001011101111101001001010000000",
		1312 => "11010111011110000111000110100111",
		1311 => "10101001011101010110111101100111",
		1310 => "01101110011001010110000101101101",
		1309 => "01110010011100100111100001110111",
		1308 => "01111001011110100111110001111110",
		1307 => "01110001100001011001100010010011",
		1306 => "10001000100110001000101001110100",
		1305 => "10001111011110100111110101111011",
		1304 => "01101101011100000111010001101111",
		1303 => "01110010011101100110101101110101",
		1302 => "01110110011101110111011101110001",
		1301 => "01110011011101010111011001101111",
		1300 => "01110010011100010110110001101110",
		1299 => "01110111011111100111111001110101",
		1298 => "01110000011010110110101001101101",
		1297 => "01101011011011000111001101110111",
		1296 => "01110110011100110111010101111010",
		1295 => "01110100011100110111000101111001",
		1294 => "01111010011101100111001001110001",
		1293 => "01111000011110000111100001110011",
		1292 => "01110001011100100111100001111001",
		1291 => "01110110011101100111010001110010",
		1290 => "01110010011100010111100001110001",
		1289 => "01110001011101100111001001111001",
		1288 => "01110100011101110111011101110111",
		1287 => "01110111011100100111011101111000",
		1286 => "01110011011101000111001001110100",
		1285 => "01110101011101110111010001110010",
		1284 => "01110100011101000111011101110010",
		1283 => "01110010011101000111001101110010",
		1282 => "01110101011100010111100101110111",
		1281 => "01110101011100010111000001110010",
		1280 => "11111110000000000000000000000000",
		1220 => "01110101011100010111001001110111",
		1219 => "01110101011100000110110101110101",
		1218 => "01110101011011110111001001110011",
		1217 => "01101111011001100111011001101110",
		1216 => "01110010011100010111011001101111",
		1215 => "01110010011011110111100001111000",
		1214 => "01110100011101000111011101110100",
		1213 => "01111000011110000111000101110110",
		1212 => "01110101011010100110011001100110",
		1211 => "01011010010101000101100101011001",
		1210 => "01010111010011100101100101100011",
		1209 => "01011110010111100101110101100100",
		1208 => "01100111011100000111010101111010",
		1207 => "01110001011101000111010001110011",
		1206 => "01110011011101000111000001110001",
		1205 => "01110001011100000110010101101010",
		1204 => "01100010011100100111001001110011",
		1203 => "10000110100000101000001001110001",
		1202 => "01110111100001100111000101100101",
		1201 => "01100111011010110111001101111000",
		1200 => "01110111011101000111100101110111",
		1199 => "01110110011101010111100101110011",
		1198 => "01110011011110000111101101111000",
		1197 => "10000011011110010111010010001000",
		1196 => "01110010100000110111011101110000",
		1195 => "10110111011100111000101101111000",
		1194 => "01111011011110010111001101110000",
		1193 => "01110100011110000111011001110010",
		1192 => "01111000011110010111010101101111",
		1191 => "01100111011010101000100110001000",
		1190 => "10001011100100110111101010001100",
		1189 => "01110001011110110111000101101110",
		1188 => "01110001011101101000001110000011",
		1187 => "01111100011111000110101001110100",
		1186 => "01110001011110010111011101110010",
		1185 => "01110010011110000110111101101111",
		1184 => "01110001100000111001010001111001",
		1183 => "10011101011101110111111001101110",
		1182 => "01101011011011000111000001101000",
		1181 => "01101111011011110110110101110010",
		1180 => "01101101011010100110011101101101",
		1179 => "01110010011110100111100101111000",
		1178 => "01110111011110000110101101101101",
		1177 => "01110111011110110111111010000111",
		1176 => "10000010011101101000010001100111",
		1175 => "01111011011011010110011101110000",
		1174 => "01110110011100110111100110001101",
		1173 => "01101000011001000111010001101110",
		1172 => "01101111011101110111000101110001",
		1171 => "01111000011101100110100101100101",
		1170 => "01100001011010110111101001110011",
		1169 => "01110001011111101000101110001111",
		1168 => "01110111011100010110010001101111",
		1167 => "01110101011010100111000101101001",
		1166 => "01101010011100100110100001111001",
		1165 => "01111100011110000111010101110110",
		1164 => "01110010011100110110100001100101",
		1163 => "01011101010110011000000001101111",
		1162 => "01110001011101010110111001110110",
		1161 => "01110101100100000110101101011110",
		1160 => "01110111011010110110101001101100",
		1159 => "01111000100011101000100101110101",
		1158 => "01111110011100000111011001110010",
		1157 => "01110010011101010101110101100010",
		1156 => "01101110011000101000011110000011",
		1155 => "01110111011100010110101010010010",
		1154 => "10000000100001101001100010100010",
		1153 => "01110101011011001000110110001010",
		1152 => "10001000100001000111110101111010",
		1151 => "01101100011110000111001001110110",
		1150 => "01101111011011100101111101100001",
		1149 => "01110011011101001001000101111100",
		1148 => "01101011100110001000111110001111",
		1147 => "10001100101001000111111101110111",
		1146 => "01111110100001111000111010010010",
		1145 => "10001111011110100111010001101011",
		1144 => "01011100011101000111100101111001",
		1143 => "01110100011010000110100101100101",
		1142 => "01111010011110011000111110011100",
		1141 => "10000011100000111001001110001111",
		1140 => "10100011100011110111111010001010",
		1139 => "01111100011111111000011110010111",
		1138 => "10010111100000100111000101011010",
		1137 => "01101001011100010111011101110110",
		1136 => "01110000011100110110010101001000",
		1135 => "01111011100110100111010101110000",
		1134 => "10010001011111111010000110100001",
		1133 => "10001001100001000110011110001000",
		1132 => "10100001100011111001100010010000",
		1131 => "10010011100100101000010010001111",
		1130 => "01111110011110100111100101110100",
		1129 => "01111000011010000111001001101000",
		1128 => "01110011100011001000010010000110",
		1127 => "10100101100000001010001010010100",
		1126 => "10000111100000010110101110101111",
		1125 => "10010011100010011000011110000110",
		1124 => "10011000100100111010001010011111",
		1123 => "01101111011011000111011001111000",
		1122 => "01101111011101000111000101100100",
		1121 => "01110100100101001010010010011011",
		1120 => "01111111100011001000101010001101",
		1119 => "10100100011101100110110010101101",
		1118 => "10100100101000011001110010001100",
		1117 => "10011010100111101000100101110101",
		1116 => "01101000011011100111010101110110",
		1115 => "01110100011010110110110001110110",
		1114 => "01101111100011101010100110001100",
		1113 => "10001000011110110111100010001111",
		1112 => "10000110011001110111011011011101",
		1111 => "10011101101001110111110010101011",
		1110 => "10110000100100101000000101011111",
		1109 => "01100011011001100111001101111000",
		1108 => "01110101011100100110001101010101",
		1107 => "01011100011101000110111001110110",
		1106 => "01111101100000001000111110100011",
		1105 => "10100101010101100100110010110110",
		1104 => "01111011101101001010101110010001",
		1103 => "10001110100011111000000001100100",
		1102 => "01101111011011000110111101111001",
		1101 => "01110100011011110110011001101010",
		1100 => "01100011100001101000101101110111",
		1099 => "10010001011111110111111101100110",
		1098 => "01101111010100010110010110010001",
		1097 => "01111100011100111000100101111001",
		1096 => "01111001011011010110011101101000",
		1095 => "01101001011011110111001001111000",
		1094 => "01110001011100100111000001101101",
		1093 => "10000111011111101000100010000111",
		1092 => "01111011100011010111100110001001",
		1091 => "01101010010111010110111101101110",
		1090 => "01111011011011100111010101111111",
		1089 => "01111010011110000111111001101000",
		1088 => "01101100011101100111011001110010",
		1087 => "01110110011100001000111010001101",
		1086 => "10001011011010001000100101110110",
		1085 => "01110000100000000111001001100111",
		1084 => "01101010011001010110100001101011",
		1083 => "01111111011011111000100001110001",
		1082 => "10001010100001111001000001111001",
		1081 => "01110101011111000111010101110010",
		1080 => "01110110011110110111101110001100",
		1079 => "10011011100011101000010001111111",
		1078 => "01111101011100110111011101100101",
		1077 => "01100111011000100110100001100011",
		1076 => "01110100011011101000001101111110",
		1075 => "10000110100001001001000110000010",
		1074 => "01110011011100100111000001110010",
		1073 => "01111001011110100111000101111101",
		1072 => "10011101100000000111001101110100",
		1071 => "01110100011010000110111001100111",
		1070 => "01100000011001110110100001101111",
		1069 => "01110010011100101000100001111101",
		1068 => "01111100011111001000110001111101",
		1067 => "01101110011100100111100001111000",
		1066 => "01110100011011100111001101111101",
		1065 => "10011001100010100111110110000011",
		1064 => "10001011100010010111111110001011",
		1063 => "01111101011111010110100110010000",
		1062 => "10000111011110111000001001111000",
		1061 => "01110100011100000111110001111110",
		1060 => "01111001011110000111001001110011",
		1059 => "01111001011100100111011010001110",
		1058 => "10010010100111111001111110011101",
		1057 => "10010011011101111000000010000010",
		1056 => "01110100011101010111110101110100",
		1055 => "01101111011000110110011001100010",
		1054 => "01110001011001100111011101111000",
		1053 => "01111001011100100111010101110111",
		1052 => "01110001011101100111100101110001",
		1051 => "01110110011101010111001101110111",
		1050 => "01110010011001100110100101100001",
		1049 => "01100000010110010011111001001110",
		1048 => "01011000010110100101010001010111",
		1047 => "01101011011011110111011101110011",
		1046 => "01110100011100110111001101110011",
		1045 => "01110001011100010111100101111000",
		1044 => "01101111011011100110111001101100",
		1043 => "01101111011010100110111001100100",
		1042 => "01100101011010100110001101011000",
		1041 => "01011110010111100110101101100110",
		1040 => "01100110011100000111100001110110",
		1039 => "01110110011110010111010001110010",
		1038 => "01111001011100100111011101111001",
		1037 => "01110101011100000111000101110011",
		1036 => "01110101011100100110111101101000",
		1035 => "01100011011101010110110101100011",
		1034 => "01101001011100100111001101101100",
		1033 => "01100111011011100111010101110110",
		1032 => "01110001011101100111100101110100",
		1031 => "01110001011101010111011101111010",
		1030 => "01110100011101000111100001111001",
		1029 => "01111000011100010111010101110001",
		1028 => "01111000011101010111000101111000",
		1027 => "01110111011110010111001101110011",
		1026 => "01110110011110010111100101111000",
		1025 => "01111001011101000111001001110011",
		1024 => "10001001000000000000000000000000",
		964 => "01110001011110010111001001110110",
		963 => "01110100011101010111101001110100",
		962 => "01110110011100100111010101110011",
		961 => "01111000011100100111000101110111",
		960 => "01110101011101000111001001110111",
		959 => "01110010011110000111100101110101",
		958 => "01111000011101100111100101111001",
		957 => "01111010011100010111000101110101",
		956 => "01111001011110010111001101111001",
		955 => "01111011100001101000100110010000",
		954 => "01111110100001001000110101111100",
		953 => "10001010011111100111010001111000",
		952 => "01110111011110010111011001110000",
		951 => "01111000011100010111011101111000",
		950 => "01110111011100010111011101110101",
		949 => "01110001011101110111001001111010",
		948 => "10100010100111001001110110101101",
		947 => "10100011100011111100100111010011",
		946 => "10101100101111001100000111001011",
		945 => "10100110100110011000000101111000",
		944 => "01101011011110100111010001111001",
		943 => "01110010011100010111001001110000",
		942 => "01110011011110001000000101111100",
		941 => "01110011011011011010000010100101",
		940 => "01111101101100011001110010000000",
		939 => "10011111100111100111111110001011",
		938 => "10011110101000101000010010011000",
		937 => "10001010011110010111100101110001",
		936 => "01111000011101010111001001101111",
		935 => "01101101011011100111010010000100",
		934 => "01111111101110010111001001101000",
		933 => "01111000011011011001000101101000",
		932 => "10010110100010111000101110000000",
		931 => "10010101100011111000110010011010",
		930 => "10010100100000010111011001110011",
		929 => "01111010011101000110111101101101",
		928 => "01110000100001110111010110011000",
		927 => "01111111011101011001010001111110",
		926 => "10001000011011100110111101101111",
		925 => "10001010011101111000001101111101",
		924 => "10001101100011000111100110000110",
		923 => "10001011011111110111010101111000",
		922 => "01110000011100100111011001100110",
		921 => "01110010100000100111000101101101",
		920 => "10101100100011110111101110000111",
		919 => "01111101011100010111010101110101",
		918 => "01110101011101100110011110001011",
		917 => "10011001100100010111000010001101",
		916 => "10001110011110000111011101110100",
		915 => "01110001011101000110111101110010",
		914 => "10001110100000011001001110111110",
		913 => "01111011100110111000101001111110",
		912 => "01110101100001100111001101100011",
		911 => "01111001011111111010110110001111",
		910 => "10010011101011101001100010011001",
		909 => "10010110011100100111001101111001",
		908 => "01110110011100110110110101110010",
		907 => "10011000011110011000110001110010",
		906 => "10001111100010101001011101111110",
		905 => "01110101011110010111110001110011",
		904 => "01110000100000110111010110000001",
		903 => "01110101011101111010000010001101",
		902 => "10010111011011010111000001111001",
		901 => "01110011011101110110110001100110",
		900 => "01111111101001101001111101111110",
		899 => "10000000011111111000001010100000",
		898 => "10001001011001110110101101101000",
		897 => "01101111011011010110100101111010",
		896 => "01111000101010001001100010001110",
		895 => "10100100011110010111001101110010",
		894 => "01110011011011110110010101101110",
		893 => "10011110100001010111111001110010",
		892 => "10100000011101101001100101110110",
		891 => "01100101011001000110011001100111",
		890 => "01101001011010000110011101110001",
		889 => "10001010011101011000010110100001",
		888 => "10010010011110100111100101110100",
		887 => "01110011011100100110100110100111",
		886 => "10100111100101101000000010001100",
		885 => "10010010100110000111110001100110",
		884 => "01110100011101001011111101110001",
		883 => "01111111011110110111101001100111",
		882 => "01101111011100101001000010010101",
		881 => "01111111011111110111010001111000",
		880 => "01110110011100100110111010010000",
		879 => "10100010100100101001000010100111",
		878 => "01111100011011100111111001111111",
		877 => "10001100100001110111001010000110",
		876 => "10000000011100100110111101101000",
		875 => "01101110011110000111000001111001",
		874 => "01111000011101010111100101110001",
		873 => "01110100011100010110111101110110",
		872 => "01110010011010010111111001101111",
		871 => "01101000100000100111111001111100",
		870 => "10000001100001011000010010010101",
		869 => "01110011011110110111101001110100",
		868 => "01101111011010110110011001101011",
		867 => "01111100011110010111011001110110",
		866 => "01110010011110010111101101110000",
		865 => "01100111010101010110100101110001",
		864 => "01111100100010110111101110001010",
		863 => "01110000100100001001111010001100",
		862 => "01111011011100100111001001110011",
		861 => "01110110011101000110111101101000",
		860 => "01110111011110010111010001110100",
		859 => "01110001011100010111100001101100",
		858 => "01100101011010000110100101111010",
		857 => "01110111100001110111011010001110",
		856 => "10000110100111110111111010010100",
		855 => "01111000101000000111001101101111",
		854 => "01111000011100010111000101110110",
		853 => "10000000011100000111000101110111",
		852 => "01110110011100000111100001100001",
		851 => "01110010100100100111000011000011",
		850 => "01111010011111101001100001110110",
		849 => "10010011100100111001011110000100",
		848 => "01110100011001110110101001110001",
		847 => "01101110011101100110111110001111",
		846 => "10011000011100100111000001110010",
		845 => "01110000011100110111001001100100",
		844 => "10000001100110110111010010001011",
		843 => "10001001100011101000100110010001",
		842 => "01110101011101111000100001100010",
		841 => "01100111011001100110011001101101",
		840 => "01110010100000010111000010001010",
		839 => "10010100011101010111000001110111",
		838 => "01110010011100100111000101011000",
		837 => "01101100101011111000000010101001",
		836 => "10001111011111111000100010010110",
		835 => "10100010100110010110100101101010",
		834 => "01100100011100111000001010001100",
		833 => "10011000100100011000101110101001",
		832 => "10000101011101010111011101110010",
		831 => "01110001011100010110111101011110",
		830 => "01100010101010001000001101111110",
		829 => "10000100100111110111111010001000",
		828 => "01111010100000101000000110000101",
		827 => "01111001100011110110110101110001",
		826 => "01111001011101010111111110010101",
		825 => "01111011011100110111010001110110",
		824 => "01110001011101010110111101110000",
		823 => "01110011011011100110100001111111",
		822 => "10001000011010101000101101111000",
		821 => "10000111100101100111000110001010",
		820 => "01110101011101111000011010010010",
		819 => "10001010100010011001101010001010",
		818 => "10000000011101010111101001110011",
		817 => "01110010011101110111010101110011",
		816 => "01111001011110111000110110000101",
		815 => "01101000101001010111000110001100",
		814 => "10000101011101101010000101110111",
		813 => "10000111100101111001011110000010",
		812 => "01111001100010011000001010000001",
		811 => "10000100011101010111010001110001",
		810 => "01110010011110000111010001101110",
		809 => "01101111011101100111010101110110",
		808 => "10011111011111000111001110100011",
		807 => "10000110011111001000100010010000",
		806 => "10010001100010101000011101111111",
		805 => "10001110100101011001101010010000",
		804 => "01111101011110010111100101110101",
		803 => "01110001011101100111001001101111",
		802 => "01100100011101000111010101110110",
		801 => "10010001101010101000100010111111",
		800 => "10011111100110101010100010101100",
		799 => "10101001101001011000111110010100",
		798 => "10001011100010111000110101111001",
		797 => "01110111011100010111010101111000",
		796 => "01110100011101000111011101110111",
		795 => "01110000011010100111000110011101",
		794 => "10010010100100111001100110011001",
		793 => "10011000101100111000110010101000",
		792 => "10011110100100001000000110001100",
		791 => "10000001100000101000010001110111",
		790 => "01110001011110010111001001110010",
		789 => "01110111011100100111010101110010",
		788 => "01110101011101010111000101111000",
		787 => "01110001011011110111000001110000",
		786 => "01101101011100100111010101111101",
		785 => "01110111011100010111010101110100",
		784 => "01110100011101100111100001110001",
		783 => "01110001011100110111100001111000",
		782 => "01110111011110000111100101110011",
		781 => "01110111011101010111001001110001",
		780 => "01110011011101110111000101110100",
		779 => "01111001011100100111001101110010",
		778 => "01110010011110010111001001110011",
		777 => "01110110011110010111001001110011",
		776 => "01110110011110100111100001111001",
		775 => "01111000011100110111011001111001",
		774 => "01110110011100110111100001110011",
		773 => "01110111011101010111001001110100",
		772 => "01111001011100110111100101110111",
		771 => "01111001011101100111011001110001",
		770 => "01110110011100100111001001110000",
		769 => "01110101011101000111000101110100",
		768 => "01010011000000000000000000000000",
		708 => "01110101011100010111100001110110",
		707 => "01110110011101100111011001110110",
		706 => "01110111011101100111010001110010",
		705 => "01110110011101000111100101111000",
		704 => "01111010011100010111011101110110",
		703 => "01110100011110000111100101111000",
		702 => "01110001011101010111010001110100",
		701 => "01111000011100010111010101110001",
		700 => "01110101011100110111001101110100",
		699 => "01110010011011010110110001101110",
		698 => "01101100011011100110111001110000",
		697 => "01110001011101000111011101101110",
		696 => "01110000011110010111000001110110",
		695 => "01111000011110000111001101110111",
		694 => "01111000011111000111011001111000",
		693 => "01110010011001010110010101100100",
		692 => "01100101011011100111111110001000",
		691 => "10010101100010110111010101110100",
		690 => "01101000011001110101110001011110",
		689 => "01101010011011110110111001110001",
		688 => "01101111011101000111011101110100",
		687 => "01110011011110001000100110010111",
		686 => "10000000100000001000111010000000",
		685 => "10000100101001101010101001110010",
		684 => "01101011111111110110010010100000",
		683 => "01110111011111111000101101111001",
		682 => "01101111011001110110000101101101",
		681 => "01101010011100100111010101110111",
		680 => "01110110011101010111111110001100",
		679 => "10010001100111001001111110010001",
		678 => "10101011101001010110111110001001",
		677 => "01101110011100100110101010001101",
		676 => "10010010011011111001011101111001",
		675 => "10010011011111110111011001111001",
		674 => "01110110011110010111000101110010",
		673 => "01110011011100011000000010000110",
		672 => "10000011100011001000000010010100",
		671 => "01111000100011010111000101111110",
		670 => "01110010011110000111101001111011",
		669 => "01111111100000001001101110100011",
		668 => "10100011100111111000010110001110",
		667 => "10000010011111110111011101110110",
		666 => "01110101011101111000011010000111",
		665 => "10011111100100111000110001111101",
		664 => "10111100100011011010010010000111",
		663 => "01101100011111111000101001110001",
		662 => "10000111100000011001100001100110",
		661 => "10000101100010111000000110000011",
		660 => "10000010100000110111100001110101",
		659 => "01110100011110011000011110010100",
		658 => "10001000100011111001110110100000",
		657 => "10011000100001100110110101111010",
		656 => "10000101011011100111101010000110",
		655 => "10101100100010101001110110010111",
		654 => "10111100100111101001011110010010",
		653 => "10000001100000000111001001110111",
		652 => "01111010100001001010100110000100",
		651 => "10001111100111111000110110000010",
		650 => "01101100100010011000111110001100",
		649 => "10001010011111011010011101111100",
		648 => "10000000101000001001101010001011",
		647 => "10001100011110001000101010001111",
		646 => "01101100011100100111011101110100",
		645 => "01110111011110101010100010101111",
		644 => "10100001100100101000100101110100",
		643 => "10001110011110011001101110000000",
		642 => "01101111100001011000001010110110",
		641 => "10000000100100110111100101111111",
		640 => "10101100100101111010111110010101",
		639 => "10000000011101110111001001110001",
		638 => "01111101100100111100100110001101",
		637 => "01110000011111110111010101111011",
		636 => "01111011011111100110011001110101",
		635 => "10010010011110011000110110001101",
		634 => "10001100101100011000110101111111",
		633 => "10010010100101001000101010010011",
		632 => "10010011100000000111001101110100",
		631 => "01111101101011111100000010100000",
		630 => "10001111101000001011101101101101",
		629 => "10001010011101001100011101111101",
		628 => "01110011100011101010000110010110",
		627 => "10001011100000001001111001101110",
		626 => "01111111100111101000010010011101",
		625 => "10011001011100110111001001111000",
		624 => "10000000100110111010011010100101",
		623 => "01101001011001110110111101101100",
		622 => "10000000011011110110101001111100",
		621 => "10000101011111101000011101111000",
		620 => "10001000011111011000000110001100",
		619 => "01111100101000011010000010001001",
		618 => "01110111011100010111011001110101",
		617 => "01111001100110001001110010010000",
		616 => "10001101011100110110111110001111",
		615 => "01110100100011010110101101111110",
		614 => "01110111100000011001000001111100",
		613 => "10001101100000100110111101110000",
		612 => "10000100011010000101010001010111",
		611 => "01101000011101010111100001110011",
		610 => "10001001101010001011000110111001",
		609 => "01111001100000011000111001101111",
		608 => "01101111011010010111011101110110",
		607 => "01101001011111001010001001111010",
		606 => "10010010011011010110101101101101",
		605 => "01011100010011010100001101000101",
		604 => "01100101011110010111011101110011",
		603 => "01110111100011101010001010000101",
		602 => "01100111011110111000111101111110",
		601 => "10010101011001010110101001110010",
		600 => "01100110011001100110100001101000",
		599 => "01100011011010000110100101101010",
		598 => "01011010010101000110010001100101",
		597 => "01100110011101100111001101111001",
		596 => "01110100011110000111110101101110",
		595 => "01110100011111101000101101110100",
		594 => "10011100011100110110001101110011",
		593 => "01101000011001000101110101100001",
		592 => "01100011010111010110101001101100",
		591 => "01110101100000001000000001101111",
		590 => "01110010011101110111010101110111",
		589 => "01111000011110100111000101011010",
		588 => "01110100011101001000000110000110",
		587 => "01110011100000001001101101111011",
		586 => "01101000011100100110110001111101",
		585 => "10000000011101010110111101111110",
		584 => "01111110101100111001101101101101",
		583 => "01111011011011110111011101111001",
		582 => "01110110011100010110100101011010",
		581 => "01111110100010110111010101111011",
		580 => "01110110100011000111101110001110",
		579 => "10010110100011110111011001111010",
		578 => "01101100100010011001010001110010",
		577 => "01110010011001011001111110001001",
		576 => "01111000011101100111000001110100",
		575 => "01110101011100100110011101011011",
		574 => "10000001011111010111001110001001",
		573 => "10100001011001111000011101110011",
		572 => "01111000011101100111000001101110",
		571 => "10000000100110110110111010000011",
		570 => "10000111011110011000000110010111",
		569 => "01111001011100110111010101110100",
		568 => "01110101011100010111001001011110",
		567 => "01011001100111011000000001101100",
		566 => "01101100011111010110010001111110",
		565 => "01101110011110111001101101101110",
		564 => "10000110011011100111010110011100",
		563 => "01110010100100011000100010011001",
		562 => "01111001011111000111011001110111",
		561 => "01110011011100010111001101100000",
		560 => "01011111011011100111001001110000",
		559 => "01110100011111010111010010000100",
		558 => "10000000011101100111110101111100",
		557 => "01110001100110011001010101110111",
		556 => "10001000011111010111101110000010",
		555 => "01110111011100100111001101110110",
		554 => "01110011011101110111001101100011",
		553 => "01101100011101100111111110001101",
		552 => "10000011100000101000010110011010",
		551 => "01111110100000001000100010001111",
		550 => "10011100011111100111101010001100",
		549 => "01111111011110000111110001110011",
		548 => "01110111011101110111100101110100",
		547 => "01110111011100010111011001100110",
		546 => "01011111011000000110110001110111",
		545 => "01111101100100101001101110100000",
		544 => "10010101101110001001000010101000",
		543 => "10100110100110001001101010000110",
		542 => "10000110100011110111010001101111",
		541 => "01110110011101100111010101110111",
		540 => "01110101011110000111001101110010",
		539 => "01101101011011100110111101101110",
		538 => "01110100011100111000100110010110",
		537 => "10000111100100001010001110001111",
		536 => "10010111100101011001110010000000",
		535 => "01111101011100100111100001111001",
		534 => "01110110011100100111000101110010",
		533 => "01111001011100100111100101111010",
		532 => "01110000011101000111010001110010",
		531 => "01101111011100101000000001111101",
		530 => "10001010011101110111101010000110",
		529 => "10000011011111111000001101110100",
		528 => "01110011011100110111011001110100",
		527 => "01110010011101110111001001110101",
		526 => "01110001011100110111010001110111",
		525 => "01110100011110000111001101110010",
		524 => "01111000011100110111001110000010",
		523 => "01111110011101100111001001101111",
		522 => "01110111011011110111011101110011",
		521 => "01110111011101100111100001110111",
		520 => "01110100011100100111011101111001",
		519 => "01111010011101010111000101111001",
		518 => "01111000011110000111101001110010",
		517 => "01111010011101110111001101110110",
		516 => "01111001011100100111001001111000",
		515 => "01110100011100010111010101110100",
		514 => "01111001011110000111100101111010",
		513 => "01110110011100100111001001110111",
		512 => "10000011000000000000000000000000",
		452 => "01110011011100010111010001110011",
		451 => "01110100011101110111011101110011",
		450 => "01110100011100000111000101110001",
		449 => "01111010011101110111000001110100",
		448 => "01111001011100010111100001110101",
		447 => "01110111011101100111001001110110",
		446 => "01110001011100010111010001110110",
		445 => "01110100011101100111011101110110",
		444 => "01110011011101000111001101110000",
		443 => "01101111011100000111001101101110",
		442 => "01110001011010010110100101101101",
		441 => "01101011011010110110111101101111",
		440 => "01110011011101100111001101110110",
		439 => "01110110011101000111100001110011",
		438 => "01110100011110010111011101111001",
		437 => "01111001011101000111100101101110",
		436 => "01101011011001100110000101011000",
		435 => "01100001011010000110110001101000",
		434 => "01011001010011010110101101101000",
		433 => "01101000011010110110011101110001",
		432 => "01110010011110000111100001110110",
		431 => "01110101011100100111100101110011",
		430 => "01110000011010110111010001110010",
		429 => "01111101011111010111100001010111",
		428 => "01110000011101000110011001101100",
		427 => "01100110011100010111100001101001",
		426 => "01110101011100110111010001101110",
		425 => "01110000011100110111001001110010",
		424 => "01110111011110110111010001110101",
		423 => "01101011011011100110011001111010",
		422 => "10000110011100101001100101111110",
		421 => "10000101011010001000001110010010",
		420 => "10000011011110001000010001111111",
		419 => "10000010100011011000110001101100",
		418 => "01101010011101110111101001110111",
		417 => "01110010011101110111011001111011",
		416 => "01110000011001011000010110011111",
		415 => "10011000101001101001010101111011",
		414 => "01111010011101110101001000111111",
		413 => "01011111011101001000010110000110",
		412 => "10001000101001101100011010000101",
		411 => "01111010011101010111001001110100",
		410 => "01111001011110010111100110001000",
		409 => "01101110011001111001011010100010",
		408 => "10001101101001010110111001110101",
		407 => "10001010100010010111110110000000",
		406 => "01111111100100001000010010001010",
		405 => "10011011101000001010001110000001",
		404 => "01111111011100100111010001110101",
		403 => "01111001011110110111110010000000",
		402 => "01110101011110101000110110010010",
		401 => "10011100101011001010011110011000",
		400 => "01101110011110000111010110000011",
		399 => "10001100100100001000101110010111",
		398 => "10001100011110000101001101110000",
		397 => "01110111011101110111100001110100",
		396 => "01110100011110010111110110001010",
		395 => "01111111011110000111010110001000",
		394 => "10010110011111100110100110011001",
		393 => "10000000011101011000011001111000",
		392 => "01111001100001111001000101111011",
		391 => "10001000011011000101001001101001",
		390 => "01110100011101010111010001110100",
		389 => "01110011011101100111101010000001",
		388 => "01111001011110001000001110001110",
		387 => "01110100011110000111000101011000",
		386 => "01100011100100011000110010000100",
		385 => "01110101011110001000010010000101",
		384 => "01101000010100010101110101110100",
		383 => "01111000011101100111010001110101",
		382 => "01111001011100100111000001111010",
		381 => "01110111011111010111010001110100",
		380 => "01101110011010110101101001100110",
		379 => "10000010100101101001000110001001",
		378 => "01110011100010110111010101110110",
		377 => "01101011010111100110011101110001",
		376 => "01110000011101010111000001111001",
		375 => "01110110011101100111000001111001",
		374 => "01101011011010100111001101101001",
		373 => "01011101010111010101011101111010",
		372 => "01110000101010011001001001110110",
		371 => "01111010011101101000010101110101",
		370 => "01101011011001100111000101111000",
		369 => "01110101011110100111100001110101",
		368 => "01110011011101110111011101110001",
		367 => "01101111011011100111000001011111",
		366 => "01010110010111100110011010100011",
		365 => "10000101101011001001010010010010",
		364 => "01111000011010000110111010000101",
		363 => "01110010011010100110110101110111",
		362 => "01110010011110010111100001110010",
		361 => "01110101011110010110111101110010",
		360 => "01101111011011110110111001101100",
		359 => "01011111011000110110111110000101",
		358 => "10010010101000111001000110001000",
		357 => "01100101010110110111000010000001",
		356 => "01101010011100110111010001110111",
		355 => "01111001011100110111000101111001",
		354 => "01110110011101010111001001101100",
		353 => "01110000011011110111010101101111",
		352 => "01101000011011101010000010000111",
		351 => "10010101101000101001010110001011",
		350 => "01100111010110110111100110001000",
		349 => "01110111011101100111100101111100",
		348 => "01110101011110000111011001111000",
		347 => "01110111011101010111010101110000",
		346 => "01110110011101110111011101110101",
		345 => "01101110011101101000000110001010",
		344 => "10011110101011011001100010000111",
		343 => "01101111011100100111110101110101",
		342 => "01111100011110000111010001110101",
		341 => "01111000011100010111100001110001",
		340 => "01110010011101100111001101100110",
		339 => "01101100011010010111000101110110",
		338 => "01110101011111100111001110010000",
		337 => "10101011101010001001110101111010",
		336 => "01110101011101110111001101110010",
		335 => "01101010010110100110101101110000",
		334 => "01110100011101110111011001110110",
		333 => "01111001011101110110110101100011",
		332 => "01100001011001110111011101101010",
		331 => "01110111011100111000100010010001",
		330 => "10101000100100111001001001111001",
		329 => "10001101011110110111001001111000",
		328 => "01101000010110010101101001100111",
		327 => "01110100011101100111100101110010",
		326 => "01111000011100010110011101100101",
		325 => "01100010011011010111001101101011",
		324 => "01101110011110011000000110001101",
		323 => "10010010100010000111101101110001",
		322 => "01110011011100110111000001110100",
		321 => "01110101011001010101100001101101",
		320 => "01111000011101100111011001111001",
		319 => "01111001011011110110011001010010",
		318 => "01011111011100010110111001101100",
		317 => "01111101011101101000011001101010",
		316 => "10000100011111000111110001111001",
		315 => "01101010011100010110011101101000",
		314 => "01101111011000100110010101110110",
		313 => "01111000011011010111001001110011",
		312 => "01110010011101100110001001011100",
		311 => "01110001011101101000000010000100",
		310 => "01111111011100000110111001111000",
		309 => "01011000011111000110100110000000",
		308 => "01101101011100100110111101100001",
		307 => "01101111011000000110011001111001",
		306 => "01110100011011110111000101110101",
		305 => "01110101011101110110010101111001",
		304 => "10000001011111100111110101111111",
		303 => "01101010100000000101101001110011",
		302 => "01100001011010100110110101110000",
		301 => "01110111011100100110101001101000",
		300 => "01100111011100010111010101110110",
		299 => "01110011011100000111011101110101",
		298 => "01110111011011110110001101101110",
		297 => "01111111100010101000100001111111",
		296 => "01111101011111010110101001111100",
		295 => "10000101011101010111101001101101",
		294 => "01101010011100010110100001100111",
		293 => "01111001100001001000000001111010",
		292 => "01111010011110000111001001110111",
		291 => "01110110011100110110100101010101",
		290 => "01101010011011010111100101111110",
		289 => "10000011011111001000001110001010",
		288 => "10000111100010101001000110000011",
		287 => "01110110011110010111001101111100",
		286 => "01110010011111100111101001110001",
		285 => "01110010011101110111100001110100",
		284 => "01110011011101010111011101110000",
		283 => "01101111011011010110101001110010",
		282 => "01110100011001110111011010001101",
		281 => "10000100011101000111110001110101",
		280 => "01100010011001100110111001110000",
		279 => "01110100011101000111100001110100",
		278 => "01110111011100000111011001110011",
		277 => "01111001011110000111100101110101",
		276 => "01111001011100110111000101111000",
		275 => "01110100011110000111011010001000",
		274 => "10010010011111111000001101110001",
		273 => "01110000011011010110111101110101",
		272 => "01110100011100100111100001110100",
		271 => "01110110011101100111100101111000",
		270 => "01111001011100100111001101110001",
		269 => "01110101011101000111000101111001",
		268 => "01111010011101010111001101110100",
		267 => "01111010011110100111011101110001",
		266 => "01111010011110000111011001110100",
		265 => "01110010011101110111010101111000",
		264 => "01110111011101000111100001110011",
		263 => "01110110011110010111010001110111",
		262 => "01110100011100010111011101110111",
		261 => "01111000011101110111000101110111",
		260 => "01111000011101110111000101110001",
		259 => "01110110011100010111000101110100",
		258 => "01110010011110010111001001110011",
		257 => "01111000011101000111010001110111",
		256 => "10111001000000000000000000000000",
		196 => "01110001011101010111100001111010",
		195 => "01110101011011010111011001110101",
		194 => "01111001011110000111011001110101",
		193 => "01110011011100010111100101110001",
		192 => "01110100011100100111011101110011",
		191 => "01110100011110010111010001111001",
		190 => "01110111011101010111100101110001",
		189 => "01110111011101000111100101111001",
		188 => "01110111011100010110110001101110",
		187 => "01110000011100010110110001101110",
		186 => "01101110011011100110101101110110",
		185 => "01110100011011100111000001101111",
		184 => "01110101011101100111011001110001",
		183 => "01110110011100010111011101110100",
		182 => "01110001011110000111100001111000",
		181 => "01110111011011010110011001100110",
		180 => "01100101010110110101101101100100",
		179 => "01011011010110110110000101011110",
		178 => "01100010010111010110011101100110",
		177 => "01101010011011000110111101110000",
		176 => "01110111011101000111011101111001",
		175 => "01110101011101100111001101110001",
		174 => "01110100011010000110010101011011",
		173 => "01100000011101001000001110000011",
		172 => "10001101100110001001101110011110",
		171 => "01110101100011001000011101111011",
		170 => "01101100011011100111001001110010",
		169 => "01110101011101000111100001110101",
		168 => "01110001011100100111010001101101",
		167 => "01101110011101000110100101100110",
		166 => "01101110011100001000111001110010",
		165 => "01111110100010011000011110000101",
		164 => "10011001100110011000111110000101",
		163 => "10001101011110000110100001100000",
		162 => "01110011011110010111011001110011",
		161 => "01110100011100010110111101101000",
		160 => "01110111100001000111011001111001",
		159 => "10000101011100111000101101111110",
		158 => "10000001011110011010100110000010",
		157 => "01110111100010101000100110001100",
		156 => "01111111100011001000000001011110",
		155 => "01110110011101010111011101110111",
		154 => "01110100011111010111001001101000",
		153 => "01101110011111110111101101111001",
		152 => "01110010011100110110111001111100",
		151 => "01111011011100000111010010010011",
		150 => "10001101100010100111110101111000",
		149 => "10010011100011001000011001110101",
		148 => "01110110011100010111011001110110",
		147 => "01110101011101000111001001101110",
		146 => "01101101100101011000100001111111",
		145 => "10000000011111101000000101101101",
		144 => "10000000011100101000100010100111",
		143 => "10010011100101111001001110010100",
		142 => "10001010100100001001010010000011",
		141 => "01101111011110010111010101110110",
		140 => "01111001011100110111000101110111",
		139 => "01111110100110011000110110000001",
		138 => "01101110100000110111111101101001",
		137 => "01101101011011000110100010011010",
		136 => "10011100100011010111101110010010",
		135 => "10010010100100111000001101111110",
		134 => "01101101011100010111011001110010",
		133 => "01110011011110000111000001111011",
		132 => "10000011100100100111010101101111",
		131 => "01110001011101010111101001110101",
		130 => "01110000011010000110000001101110",
		129 => "01111010101001111001011110011001",
		128 => "10000101100011000111111110000001",
		127 => "01110000011101010111100101111000",
		126 => "01110101011100010110111101111101",
		125 => "10000011100010110111100110001101",
		124 => "10000000011101001001110101110010",
		123 => "01101000011000100101111001110100",
		122 => "10000010101100001001011101111001",
		121 => "10001111100110011001000110000101",
		120 => "01110101011101000111100101110010",
		119 => "01110010011101000110101110000010",
		118 => "10001000100011001000100110010001",
		117 => "10000000100000101000001001101011",
		116 => "01101010010111000101100001101011",
		115 => "10010111100011001001000110011001",
		114 => "10001111100100001001010010001000",
		113 => "01110010011100110111100001110100",
		112 => "01110110011100000111110010011001",
		111 => "10010010100010001000001110010001",
		110 => "01110011011111100111000001100010",
		109 => "01011010010011100110010001110011",
		108 => "01101100100111111001000010010010",
		107 => "10011101011101001001100110001010",
		106 => "01100111011100000111100101110110",
		105 => "01111001011101111000010010100000",
		104 => "10011000100000111000111010000111",
		103 => "01110100011110000111000101011001",
		102 => "01011001010110000110110110101111",
		101 => "10011110011011101000111010000110",
		100 => "10100001100010001001001001110000",
		99 => "01101010011100100111011101110110",
		98 => "01110110011100011000000110011011",
		97 => "10010111100011010111110101101001",
		96 => "01111001011110010110111001011011",
		95 => "01010011010110010110011010000010",
		94 => "01111010100111010111111110001001",
		93 => "10010110100111010111100110000100",
		92 => "01110101011100110111101001110001",
		91 => "01111000011011100111000110101110",
		90 => "10010011100101001001000110010000",
		89 => "10001101011101000111001101011110",
		88 => "01011001011000011000011010101000",
		87 => "10000100100000110111111001111111",
		86 => "10001110101000010111011101110000",
		85 => "01110100011101000111010001111001",
		84 => "01110100011001110110011110010010",
		83 => "10001101100101001010000110001111",
		82 => "10000010011010010111001101011100",
		81 => "01011011011011001000001001101000",
		80 => "10001000011111110111001010001111",
		79 => "10010000100001110110111001101101",
		78 => "01110101011101100111001101111000",
		77 => "01110110011001010110000110100000",
		76 => "10011000100101001000100110001110",
		75 => "01110011100101101011011001111111",
		74 => "01101110100011111000110101111001",
		73 => "10001101011100111001001001111001",
		72 => "01111100011110011000011101110011",
		71 => "01111001011101110111000101110010",
		70 => "01110010011001110101111110100011",
		69 => "10011011011100110111011110001110",
		68 => "10011001100100111001000010001000",
		67 => "01100010011101011001111101110010",
		66 => "01110010100100100111110101110000",
		65 => "01110101011100010111011101110001",
		64 => "01111110011100100111100101110011",
		63 => "01110111011001100101011010001111",
		62 => "10101000100011001001000010010000",
		61 => "01110111100001111000111110101100",
		60 => "10001101100011100110111010001100",
		59 => "01110100011110101000111110000001",
		58 => "01111010011110100111010101101100",
		57 => "01110111011100010111010101111001",
		56 => "01110001011001000101110101110001",
		55 => "10010001011100110111110001111000",
		54 => "10001000100100101001010101110000",
		53 => "01110011011111001000011001110100",
		52 => "10001000100000101000100001110000",
		51 => "10000111100000110111011101110001",
		50 => "01110100011110000111001001110011",
		49 => "01110110011011000101110001011110",
		48 => "01110011100111111001100110001000",
		47 => "01111101100011101000000010001101",
		46 => "01110010100011111001000001101111",
		45 => "01110111011111000110100001111111",
		44 => "01111110100000010111000001101111",
		43 => "01111000011101110111001101110110",
		42 => "01110010011100000110011101100110",
		41 => "01101100011110101000000001110010",
		40 => "10001001100101011001001110000101",
		39 => "10000001100100001001000101110100",
		38 => "10010011100110011000010010000001",
		37 => "01111011011101010110010101110101",
		36 => "01110101011101100111011101110111",
		35 => "01111001011101000111000101101100",
		34 => "01110101011110100111010001111001",
		33 => "10000001100010111001011110000111",
		32 => "10011000100001011001011010001001",
		31 => "10100000011111111000011001111000",
		30 => "01110110011001110110101001110010",
		29 => "01110111011100010111100001110001",
		28 => "01110001011101000111011101110100",
		27 => "01110011011011010110100101110010",
		26 => "01110010011101101000101010001111",
		25 => "10000011100100011000111101111010",
		24 => "01111100011110110111010001110101",
		23 => "01100111011011010110111001111001",
		22 => "01111000011100100111011101110010",
		21 => "01110001011101010111010101111001",
		20 => "01110011011100100111000101101110",
		19 => "01110001011100000110110101101100",
		18 => "01100111011010110110111001110110",
		17 => "01110011011100100111010101110101",
		16 => "01110101011100010111100001111000",
		15 => "01111001011101010111100001110010",
		14 => "01110010011110010111010001110101",
		13 => "01110001011100010111011101110111",
		12 => "01111000011110010111101001111100",
		11 => "01110100011100000111100001111001",
		10 => "01110101011100010111011101111001",
		9 => "01110110011101100111001101110010",
		8 => "01111000011101110111010101110110",
		7 => "01110101011101100111100101110010",
		6 => "01111001011100010111010101110111",
		5 => "01110001011110010111100001110110",
		4 => "01110101011100110111011001110101",
		3 => "01110100011110000111001101110010",
		2 => "01111000011101010111011001110001",
		1 => "01110110011101000111001001111000",
		0 => "01010000000000000000000000000000", 
        -- here ends the generated array allocation

        others => "00000000000000000000000000000000"
    );

    signal rom_index: std_logic_vector (11 downto 0);
begin
    rom_index <= (in_rom_neuron_index & in_rom_input_index); -- combine the neuron and input index to adress the array
    out_data_rom <= rom_arr(to_integer(unsigned(rom_index)));
end RTL;
