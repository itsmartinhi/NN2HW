LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
ENTITY AND2 IS
  PORT (
    x, y : IN STD_LOGIC;
    z : OUT STD_LOGIC);
END AND2;
ARCHITECTURE DATAFLOW OF AND2 IS
BEGIN
  z <= x AND y AFTER 3 ns;
END ARCHITECTURE;