LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
ENTITY XOR2 IS
  PORT (
    x, y : IN STD_LOGIC;
    z : OUT STD_LOGIC);
END XOR2;
ARCHITECTURE DATAFLOW OF XOR2 IS
BEGIN
  z <= x XOR y AFTER 2 ns;
END ARCHITECTURE;